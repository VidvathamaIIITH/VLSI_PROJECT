magic
tech scmos
timestamp 1731794669
<< nwell >>
rect -765 531 -703 558
rect -669 526 -642 588
rect -765 480 -703 507
rect -772 354 -718 416
rect -710 284 -683 346
rect -118 291 -56 318
rect -22 286 5 348
rect 69 270 96 332
rect -118 240 -56 267
rect 134 173 161 375
rect 243 301 297 363
rect 183 176 210 238
rect 305 231 332 293
rect 45 -58 107 -31
rect 141 -63 168 -1
rect 1272 -3 1334 24
rect 1368 -8 1395 54
rect 1272 -54 1334 -27
rect 45 -109 107 -82
rect 38 -235 92 -173
rect 100 -305 127 -243
rect 616 -273 670 -211
rect 678 -343 705 -281
rect 913 -355 940 -153
rect 962 -352 989 -290
rect 65 -851 127 -824
rect 161 -856 188 -794
rect 65 -902 127 -875
rect 659 -909 713 -847
rect 58 -1028 112 -966
rect 721 -979 748 -917
rect 997 -918 1051 -856
rect 1377 -907 1431 -845
rect 2219 -860 2246 -658
rect 2268 -857 2295 -795
rect 2713 -843 2740 -641
rect 3552 -680 3614 -653
rect 3648 -685 3675 -623
rect 3552 -731 3614 -704
rect 2762 -840 2789 -778
rect 1059 -988 1086 -926
rect 1439 -977 1466 -915
rect 120 -1098 147 -1036
rect 50 -1975 112 -1948
rect 146 -1980 173 -1918
rect 793 -1970 847 -1908
rect 1261 -1961 1315 -1899
rect 1663 -1958 1717 -1896
rect 2164 -1923 2218 -1861
rect 2769 -1923 2823 -1861
rect 3374 -1923 3428 -1861
rect 50 -2026 112 -1999
rect 855 -2040 882 -1978
rect 1323 -2031 1350 -1969
rect 1725 -2028 1752 -1966
rect 2226 -1993 2253 -1931
rect 2831 -1993 2858 -1931
rect 3436 -1993 3463 -1931
rect 4002 -1967 4029 -1765
rect 4051 -1964 4078 -1902
rect 4456 -1996 4483 -1794
rect 4505 -1993 4532 -1931
rect 4921 -1961 4948 -1759
rect 5878 -1775 5940 -1748
rect 5974 -1780 6001 -1718
rect 5878 -1826 5940 -1799
rect 4970 -1958 4997 -1896
rect 43 -2152 97 -2090
rect 105 -2222 132 -2160
rect 50 -3394 112 -3367
rect 146 -3399 173 -3337
rect 884 -3396 938 -3334
rect 50 -3445 112 -3418
rect 946 -3466 973 -3404
rect 1222 -3405 1276 -3343
rect 1602 -3394 1656 -3332
rect 2711 -3365 2765 -3303
rect 1284 -3475 1311 -3413
rect 1664 -3464 1691 -3402
rect 2773 -3435 2800 -3373
rect 3049 -3374 3103 -3312
rect 3429 -3363 3483 -3301
rect 4204 -3348 4258 -3286
rect 3111 -3444 3138 -3382
rect 3491 -3433 3518 -3371
rect 4266 -3418 4293 -3356
rect 4526 -3362 4580 -3300
rect 4588 -3432 4615 -3370
rect 4864 -3371 4918 -3309
rect 5244 -3360 5298 -3298
rect 6057 -3324 6084 -3122
rect 6106 -3321 6133 -3259
rect 6488 -3318 6515 -3116
rect 6537 -3315 6564 -3253
rect 6942 -3347 6969 -3145
rect 6991 -3344 7018 -3282
rect 7407 -3312 7434 -3110
rect 8552 -3190 8614 -3163
rect 8648 -3195 8675 -3133
rect 8552 -3241 8614 -3214
rect 7456 -3309 7483 -3247
rect 4926 -3441 4953 -3379
rect 5306 -3430 5333 -3368
rect 43 -3571 97 -3509
rect 105 -3641 132 -3579
<< ntransistor >>
rect -795 543 -775 545
rect -692 531 -690 551
rect -692 498 -690 518
rect -656 496 -654 516
rect -795 492 -775 494
rect -740 288 -738 328
rect -148 303 -128 305
rect -45 291 -43 311
rect -740 223 -738 263
rect -697 254 -695 274
rect -45 258 -43 278
rect -9 256 -7 276
rect -148 252 -128 254
rect 82 240 84 260
rect 275 235 277 275
rect 275 170 277 210
rect 318 201 320 221
rect 132 136 134 156
rect 165 136 167 156
rect 196 146 198 166
rect 1242 9 1262 11
rect 1345 -3 1347 17
rect 15 -46 35 -44
rect 118 -58 120 -38
rect 1345 -36 1347 -16
rect 1381 -38 1383 -18
rect 1242 -42 1262 -40
rect 118 -91 120 -71
rect 154 -93 156 -73
rect 15 -97 35 -95
rect 70 -301 72 -261
rect 70 -366 72 -326
rect 113 -335 115 -315
rect 648 -339 650 -299
rect 648 -404 650 -364
rect 691 -373 693 -353
rect 911 -392 913 -372
rect 944 -392 946 -372
rect 975 -382 977 -362
rect 3522 -668 3542 -666
rect 3625 -680 3627 -660
rect 3625 -713 3627 -693
rect 3661 -715 3663 -695
rect 3522 -719 3542 -717
rect 35 -839 55 -837
rect 138 -851 140 -831
rect 138 -884 140 -864
rect 174 -886 176 -866
rect 35 -890 55 -888
rect 2217 -897 2219 -877
rect 2250 -897 2252 -877
rect 2281 -887 2283 -867
rect 2711 -880 2713 -860
rect 2744 -880 2746 -860
rect 2775 -870 2777 -850
rect 691 -975 693 -935
rect 1029 -984 1031 -944
rect 90 -1094 92 -1054
rect 691 -1040 693 -1000
rect 734 -1009 736 -989
rect 1409 -973 1411 -933
rect 1029 -1049 1031 -1009
rect 1072 -1018 1074 -998
rect 1409 -1038 1411 -998
rect 1452 -1007 1454 -987
rect 90 -1159 92 -1119
rect 133 -1128 135 -1108
rect 5848 -1763 5868 -1761
rect 20 -1963 40 -1961
rect 123 -1975 125 -1955
rect 123 -2008 125 -1988
rect 159 -2010 161 -1990
rect 20 -2014 40 -2012
rect 825 -2036 827 -1996
rect 1293 -2027 1295 -1987
rect 1695 -2024 1697 -1984
rect 2196 -1989 2198 -1949
rect 2801 -1989 2803 -1949
rect 825 -2101 827 -2061
rect 868 -2070 870 -2050
rect 1293 -2092 1295 -2052
rect 1336 -2061 1338 -2041
rect 1695 -2089 1697 -2049
rect 1738 -2058 1740 -2038
rect 2196 -2054 2198 -2014
rect 2239 -2023 2241 -2003
rect 3406 -1989 3408 -1949
rect 2801 -2054 2803 -2014
rect 2844 -2023 2846 -2003
rect 5951 -1775 5953 -1755
rect 5951 -1808 5953 -1788
rect 5987 -1810 5989 -1790
rect 5848 -1814 5868 -1812
rect 3406 -2054 3408 -2014
rect 3449 -2023 3451 -2003
rect 4000 -2004 4002 -1984
rect 4033 -2004 4035 -1984
rect 4064 -1994 4066 -1974
rect 4919 -1998 4921 -1978
rect 4952 -1998 4954 -1978
rect 4983 -1988 4985 -1968
rect 4454 -2033 4456 -2013
rect 4487 -2033 4489 -2013
rect 4518 -2023 4520 -2003
rect 75 -2218 77 -2178
rect 75 -2283 77 -2243
rect 118 -2252 120 -2232
rect 20 -3382 40 -3380
rect 123 -3394 125 -3374
rect 123 -3427 125 -3407
rect 159 -3429 161 -3409
rect 20 -3433 40 -3431
rect 916 -3462 918 -3422
rect 1254 -3471 1256 -3431
rect 916 -3527 918 -3487
rect 959 -3496 961 -3476
rect 1634 -3460 1636 -3420
rect 2743 -3431 2745 -3391
rect 3081 -3440 3083 -3400
rect 1254 -3536 1256 -3496
rect 1297 -3505 1299 -3485
rect 1634 -3525 1636 -3485
rect 1677 -3494 1679 -3474
rect 2743 -3496 2745 -3456
rect 2786 -3465 2788 -3445
rect 3461 -3429 3463 -3389
rect 4236 -3414 4238 -3374
rect 4558 -3428 4560 -3388
rect 3081 -3505 3083 -3465
rect 3124 -3474 3126 -3454
rect 3461 -3494 3463 -3454
rect 3504 -3463 3506 -3443
rect 4236 -3479 4238 -3439
rect 4279 -3448 4281 -3428
rect 4896 -3437 4898 -3397
rect 4558 -3493 4560 -3453
rect 4601 -3462 4603 -3442
rect 6055 -3361 6057 -3341
rect 6088 -3361 6090 -3341
rect 6119 -3351 6121 -3331
rect 8522 -3178 8542 -3176
rect 8625 -3190 8627 -3170
rect 6486 -3355 6488 -3335
rect 6519 -3355 6521 -3335
rect 6550 -3345 6552 -3325
rect 8625 -3223 8627 -3203
rect 8661 -3225 8663 -3205
rect 8522 -3229 8542 -3227
rect 7405 -3349 7407 -3329
rect 7438 -3349 7440 -3329
rect 7469 -3339 7471 -3319
rect 5276 -3426 5278 -3386
rect 6940 -3384 6942 -3364
rect 6973 -3384 6975 -3364
rect 7004 -3374 7006 -3354
rect 4896 -3502 4898 -3462
rect 4939 -3471 4941 -3451
rect 5276 -3491 5278 -3451
rect 5319 -3460 5321 -3440
rect 75 -3637 77 -3597
rect 75 -3702 77 -3662
rect 118 -3671 120 -3651
<< ptransistor >>
rect -757 543 -717 545
rect -656 534 -654 574
rect -757 492 -717 494
rect -759 362 -757 402
rect -732 362 -730 402
rect -697 292 -695 332
rect -110 303 -70 305
rect -9 294 -7 334
rect 82 278 84 318
rect 147 281 149 361
rect 256 309 258 349
rect 283 309 285 349
rect -110 252 -70 254
rect 147 181 149 261
rect 196 184 198 224
rect 318 239 320 279
rect 1280 9 1320 11
rect 1381 0 1383 40
rect 53 -46 93 -44
rect 154 -55 156 -15
rect 1280 -42 1320 -40
rect 53 -97 93 -95
rect 51 -227 53 -187
rect 78 -227 80 -187
rect 113 -297 115 -257
rect 629 -265 631 -225
rect 656 -265 658 -225
rect 926 -247 928 -167
rect 691 -335 693 -295
rect 926 -347 928 -267
rect 975 -344 977 -304
rect 2232 -752 2234 -672
rect 2726 -735 2728 -655
rect 3560 -668 3600 -666
rect 3661 -677 3663 -637
rect 3560 -719 3600 -717
rect 73 -839 113 -837
rect 174 -848 176 -808
rect 2232 -852 2234 -772
rect 73 -890 113 -888
rect 672 -901 674 -861
rect 699 -901 701 -861
rect 1010 -910 1012 -870
rect 1037 -910 1039 -870
rect 1390 -899 1392 -859
rect 1417 -899 1419 -859
rect 2281 -849 2283 -809
rect 2726 -835 2728 -755
rect 2775 -832 2777 -792
rect 71 -1020 73 -980
rect 98 -1020 100 -980
rect 734 -971 736 -931
rect 1072 -980 1074 -940
rect 1452 -969 1454 -929
rect 133 -1090 135 -1050
rect 5886 -1763 5926 -1761
rect 4015 -1859 4017 -1779
rect 58 -1963 98 -1961
rect 159 -1972 161 -1932
rect 806 -1962 808 -1922
rect 833 -1962 835 -1922
rect 1274 -1953 1276 -1913
rect 1301 -1953 1303 -1913
rect 1676 -1950 1678 -1910
rect 1703 -1950 1705 -1910
rect 2177 -1915 2179 -1875
rect 2204 -1915 2206 -1875
rect 2782 -1915 2784 -1875
rect 2809 -1915 2811 -1875
rect 3387 -1915 3389 -1875
rect 3414 -1915 3416 -1875
rect 58 -2014 98 -2012
rect 868 -2032 870 -1992
rect 1336 -2023 1338 -1983
rect 1738 -2020 1740 -1980
rect 2239 -1985 2241 -1945
rect 2844 -1985 2846 -1945
rect 3449 -1985 3451 -1945
rect 4015 -1959 4017 -1879
rect 4469 -1888 4471 -1808
rect 4934 -1853 4936 -1773
rect 5987 -1772 5989 -1732
rect 5886 -1814 5926 -1812
rect 4064 -1956 4066 -1916
rect 4469 -1988 4471 -1908
rect 4518 -1985 4520 -1945
rect 4934 -1953 4936 -1873
rect 4983 -1950 4985 -1910
rect 56 -2144 58 -2104
rect 83 -2144 85 -2104
rect 118 -2214 120 -2174
rect 6070 -3216 6072 -3136
rect 6501 -3210 6503 -3130
rect 58 -3382 98 -3380
rect 159 -3391 161 -3351
rect 897 -3388 899 -3348
rect 924 -3388 926 -3348
rect 1235 -3397 1237 -3357
rect 1262 -3397 1264 -3357
rect 1615 -3386 1617 -3346
rect 1642 -3386 1644 -3346
rect 2724 -3357 2726 -3317
rect 2751 -3357 2753 -3317
rect 58 -3433 98 -3431
rect 959 -3458 961 -3418
rect 56 -3563 58 -3523
rect 83 -3563 85 -3523
rect 3062 -3366 3064 -3326
rect 3089 -3366 3091 -3326
rect 3442 -3355 3444 -3315
rect 3469 -3355 3471 -3315
rect 4217 -3340 4219 -3300
rect 4244 -3340 4246 -3300
rect 1297 -3467 1299 -3427
rect 1677 -3456 1679 -3416
rect 2786 -3427 2788 -3387
rect 3124 -3436 3126 -3396
rect 4539 -3354 4541 -3314
rect 4566 -3354 4568 -3314
rect 3504 -3425 3506 -3385
rect 4279 -3410 4281 -3370
rect 4877 -3363 4879 -3323
rect 4904 -3363 4906 -3323
rect 5257 -3352 5259 -3312
rect 5284 -3352 5286 -3312
rect 6070 -3316 6072 -3236
rect 6119 -3313 6121 -3273
rect 6501 -3310 6503 -3230
rect 4601 -3424 4603 -3384
rect 6955 -3239 6957 -3159
rect 7420 -3204 7422 -3124
rect 8560 -3178 8600 -3176
rect 8661 -3187 8663 -3147
rect 6550 -3307 6552 -3267
rect 6955 -3339 6957 -3259
rect 7004 -3336 7006 -3296
rect 7420 -3304 7422 -3224
rect 8560 -3229 8600 -3227
rect 7469 -3301 7471 -3261
rect 4939 -3433 4941 -3393
rect 5319 -3422 5321 -3382
rect 118 -3633 120 -3593
<< ndiffusion >>
rect -795 545 -775 546
rect -795 542 -775 543
rect -693 531 -692 551
rect -690 531 -689 551
rect -795 494 -775 495
rect -693 498 -692 518
rect -690 498 -689 518
rect -657 496 -656 516
rect -654 496 -653 516
rect -795 491 -775 492
rect -741 288 -740 328
rect -738 288 -737 328
rect -148 305 -128 306
rect -148 302 -128 303
rect -46 291 -45 311
rect -43 291 -42 311
rect -741 223 -740 263
rect -738 223 -737 263
rect -698 254 -697 274
rect -695 254 -694 274
rect -148 254 -128 255
rect -46 258 -45 278
rect -43 258 -42 278
rect -10 256 -9 276
rect -7 256 -6 276
rect -148 251 -128 252
rect 81 240 82 260
rect 84 240 85 260
rect 274 235 275 275
rect 277 235 278 275
rect 274 170 275 210
rect 277 170 278 210
rect 317 201 318 221
rect 320 201 321 221
rect 131 136 132 156
rect 134 136 135 156
rect 164 136 165 156
rect 167 136 168 156
rect 195 146 196 166
rect 198 146 199 166
rect 1242 11 1262 12
rect 1242 8 1262 9
rect 1344 -3 1345 17
rect 1347 -3 1348 17
rect 15 -44 35 -43
rect 15 -47 35 -46
rect 117 -58 118 -38
rect 120 -58 121 -38
rect 1242 -40 1262 -39
rect 1344 -36 1345 -16
rect 1347 -36 1348 -16
rect 1380 -38 1381 -18
rect 1383 -38 1384 -18
rect 1242 -43 1262 -42
rect 15 -95 35 -94
rect 117 -91 118 -71
rect 120 -91 121 -71
rect 153 -93 154 -73
rect 156 -93 157 -73
rect 15 -98 35 -97
rect 69 -301 70 -261
rect 72 -301 73 -261
rect 69 -366 70 -326
rect 72 -366 73 -326
rect 112 -335 113 -315
rect 115 -335 116 -315
rect 647 -339 648 -299
rect 650 -339 651 -299
rect 647 -404 648 -364
rect 650 -404 651 -364
rect 690 -373 691 -353
rect 693 -373 694 -353
rect 910 -392 911 -372
rect 913 -392 914 -372
rect 943 -392 944 -372
rect 946 -392 947 -372
rect 974 -382 975 -362
rect 977 -382 978 -362
rect 3522 -666 3542 -665
rect 3522 -669 3542 -668
rect 3624 -680 3625 -660
rect 3627 -680 3628 -660
rect 3522 -717 3542 -716
rect 3624 -713 3625 -693
rect 3627 -713 3628 -693
rect 3660 -715 3661 -695
rect 3663 -715 3664 -695
rect 3522 -720 3542 -719
rect 35 -837 55 -836
rect 35 -840 55 -839
rect 137 -851 138 -831
rect 140 -851 141 -831
rect 35 -888 55 -887
rect 137 -884 138 -864
rect 140 -884 141 -864
rect 173 -886 174 -866
rect 176 -886 177 -866
rect 35 -891 55 -890
rect 2216 -897 2217 -877
rect 2219 -897 2220 -877
rect 2249 -897 2250 -877
rect 2252 -897 2253 -877
rect 2280 -887 2281 -867
rect 2283 -887 2284 -867
rect 2710 -880 2711 -860
rect 2713 -880 2714 -860
rect 2743 -880 2744 -860
rect 2746 -880 2747 -860
rect 2774 -870 2775 -850
rect 2777 -870 2778 -850
rect 690 -975 691 -935
rect 693 -975 694 -935
rect 1028 -984 1029 -944
rect 1031 -984 1032 -944
rect 89 -1094 90 -1054
rect 92 -1094 93 -1054
rect 690 -1040 691 -1000
rect 693 -1040 694 -1000
rect 733 -1009 734 -989
rect 736 -1009 737 -989
rect 1408 -973 1409 -933
rect 1411 -973 1412 -933
rect 1028 -1049 1029 -1009
rect 1031 -1049 1032 -1009
rect 1071 -1018 1072 -998
rect 1074 -1018 1075 -998
rect 1408 -1038 1409 -998
rect 1411 -1038 1412 -998
rect 1451 -1007 1452 -987
rect 1454 -1007 1455 -987
rect 89 -1159 90 -1119
rect 92 -1159 93 -1119
rect 132 -1128 133 -1108
rect 135 -1128 136 -1108
rect 5848 -1761 5868 -1760
rect 5848 -1764 5868 -1763
rect 20 -1961 40 -1960
rect 20 -1964 40 -1963
rect 122 -1975 123 -1955
rect 125 -1975 126 -1955
rect 20 -2012 40 -2011
rect 122 -2008 123 -1988
rect 125 -2008 126 -1988
rect 158 -2010 159 -1990
rect 161 -2010 162 -1990
rect 20 -2015 40 -2014
rect 824 -2036 825 -1996
rect 827 -2036 828 -1996
rect 1292 -2027 1293 -1987
rect 1295 -2027 1296 -1987
rect 1694 -2024 1695 -1984
rect 1697 -2024 1698 -1984
rect 2195 -1989 2196 -1949
rect 2198 -1989 2199 -1949
rect 2800 -1989 2801 -1949
rect 2803 -1989 2804 -1949
rect 824 -2101 825 -2061
rect 827 -2101 828 -2061
rect 867 -2070 868 -2050
rect 870 -2070 871 -2050
rect 1292 -2092 1293 -2052
rect 1295 -2092 1296 -2052
rect 1335 -2061 1336 -2041
rect 1338 -2061 1339 -2041
rect 1694 -2089 1695 -2049
rect 1697 -2089 1698 -2049
rect 1737 -2058 1738 -2038
rect 1740 -2058 1741 -2038
rect 2195 -2054 2196 -2014
rect 2198 -2054 2199 -2014
rect 2238 -2023 2239 -2003
rect 2241 -2023 2242 -2003
rect 3405 -1989 3406 -1949
rect 3408 -1989 3409 -1949
rect 2800 -2054 2801 -2014
rect 2803 -2054 2804 -2014
rect 2843 -2023 2844 -2003
rect 2846 -2023 2847 -2003
rect 5950 -1775 5951 -1755
rect 5953 -1775 5954 -1755
rect 5848 -1812 5868 -1811
rect 5950 -1808 5951 -1788
rect 5953 -1808 5954 -1788
rect 5986 -1810 5987 -1790
rect 5989 -1810 5990 -1790
rect 5848 -1815 5868 -1814
rect 3405 -2054 3406 -2014
rect 3408 -2054 3409 -2014
rect 3448 -2023 3449 -2003
rect 3451 -2023 3452 -2003
rect 3999 -2004 4000 -1984
rect 4002 -2004 4003 -1984
rect 4032 -2004 4033 -1984
rect 4035 -2004 4036 -1984
rect 4063 -1994 4064 -1974
rect 4066 -1994 4067 -1974
rect 4918 -1998 4919 -1978
rect 4921 -1998 4922 -1978
rect 4951 -1998 4952 -1978
rect 4954 -1998 4955 -1978
rect 4982 -1988 4983 -1968
rect 4985 -1988 4986 -1968
rect 4453 -2033 4454 -2013
rect 4456 -2033 4457 -2013
rect 4486 -2033 4487 -2013
rect 4489 -2033 4490 -2013
rect 4517 -2023 4518 -2003
rect 4520 -2023 4521 -2003
rect 74 -2218 75 -2178
rect 77 -2218 78 -2178
rect 74 -2283 75 -2243
rect 77 -2283 78 -2243
rect 117 -2252 118 -2232
rect 120 -2252 121 -2232
rect 20 -3380 40 -3379
rect 20 -3383 40 -3382
rect 122 -3394 123 -3374
rect 125 -3394 126 -3374
rect 20 -3431 40 -3430
rect 122 -3427 123 -3407
rect 125 -3427 126 -3407
rect 158 -3429 159 -3409
rect 161 -3429 162 -3409
rect 20 -3434 40 -3433
rect 915 -3462 916 -3422
rect 918 -3462 919 -3422
rect 1253 -3471 1254 -3431
rect 1256 -3471 1257 -3431
rect 915 -3527 916 -3487
rect 918 -3527 919 -3487
rect 958 -3496 959 -3476
rect 961 -3496 962 -3476
rect 1633 -3460 1634 -3420
rect 1636 -3460 1637 -3420
rect 2742 -3431 2743 -3391
rect 2745 -3431 2746 -3391
rect 3080 -3440 3081 -3400
rect 3083 -3440 3084 -3400
rect 1253 -3536 1254 -3496
rect 1256 -3536 1257 -3496
rect 1296 -3505 1297 -3485
rect 1299 -3505 1300 -3485
rect 1633 -3525 1634 -3485
rect 1636 -3525 1637 -3485
rect 1676 -3494 1677 -3474
rect 1679 -3494 1680 -3474
rect 2742 -3496 2743 -3456
rect 2745 -3496 2746 -3456
rect 2785 -3465 2786 -3445
rect 2788 -3465 2789 -3445
rect 3460 -3429 3461 -3389
rect 3463 -3429 3464 -3389
rect 4235 -3414 4236 -3374
rect 4238 -3414 4239 -3374
rect 4557 -3428 4558 -3388
rect 4560 -3428 4561 -3388
rect 3080 -3505 3081 -3465
rect 3083 -3505 3084 -3465
rect 3123 -3474 3124 -3454
rect 3126 -3474 3127 -3454
rect 3460 -3494 3461 -3454
rect 3463 -3494 3464 -3454
rect 3503 -3463 3504 -3443
rect 3506 -3463 3507 -3443
rect 4235 -3479 4236 -3439
rect 4238 -3479 4239 -3439
rect 4278 -3448 4279 -3428
rect 4281 -3448 4282 -3428
rect 4895 -3437 4896 -3397
rect 4898 -3437 4899 -3397
rect 4557 -3493 4558 -3453
rect 4560 -3493 4561 -3453
rect 4600 -3462 4601 -3442
rect 4603 -3462 4604 -3442
rect 6054 -3361 6055 -3341
rect 6057 -3361 6058 -3341
rect 6087 -3361 6088 -3341
rect 6090 -3361 6091 -3341
rect 6118 -3351 6119 -3331
rect 6121 -3351 6122 -3331
rect 8522 -3176 8542 -3175
rect 8522 -3179 8542 -3178
rect 8624 -3190 8625 -3170
rect 8627 -3190 8628 -3170
rect 6485 -3355 6486 -3335
rect 6488 -3355 6489 -3335
rect 6518 -3355 6519 -3335
rect 6521 -3355 6522 -3335
rect 6549 -3345 6550 -3325
rect 6552 -3345 6553 -3325
rect 8522 -3227 8542 -3226
rect 8624 -3223 8625 -3203
rect 8627 -3223 8628 -3203
rect 8660 -3225 8661 -3205
rect 8663 -3225 8664 -3205
rect 8522 -3230 8542 -3229
rect 7404 -3349 7405 -3329
rect 7407 -3349 7408 -3329
rect 7437 -3349 7438 -3329
rect 7440 -3349 7441 -3329
rect 7468 -3339 7469 -3319
rect 7471 -3339 7472 -3319
rect 5275 -3426 5276 -3386
rect 5278 -3426 5279 -3386
rect 6939 -3384 6940 -3364
rect 6942 -3384 6943 -3364
rect 6972 -3384 6973 -3364
rect 6975 -3384 6976 -3364
rect 7003 -3374 7004 -3354
rect 7006 -3374 7007 -3354
rect 4895 -3502 4896 -3462
rect 4898 -3502 4899 -3462
rect 4938 -3471 4939 -3451
rect 4941 -3471 4942 -3451
rect 5275 -3491 5276 -3451
rect 5278 -3491 5279 -3451
rect 5318 -3460 5319 -3440
rect 5321 -3460 5322 -3440
rect 74 -3637 75 -3597
rect 77 -3637 78 -3597
rect 74 -3702 75 -3662
rect 77 -3702 78 -3662
rect 117 -3671 118 -3651
rect 120 -3671 121 -3651
<< pdiffusion >>
rect -757 545 -717 546
rect -757 542 -717 543
rect -657 534 -656 574
rect -654 534 -653 574
rect -757 494 -717 495
rect -757 491 -717 492
rect -760 362 -759 402
rect -757 362 -756 402
rect -733 362 -732 402
rect -730 362 -729 402
rect -698 292 -697 332
rect -695 292 -694 332
rect -110 305 -70 306
rect -110 302 -70 303
rect -10 294 -9 334
rect -7 294 -6 334
rect 81 278 82 318
rect 84 278 85 318
rect 146 281 147 361
rect 149 281 150 361
rect 255 309 256 349
rect 258 309 259 349
rect 282 309 283 349
rect 285 309 286 349
rect -110 254 -70 255
rect -110 251 -70 252
rect 146 181 147 261
rect 149 181 150 261
rect 195 184 196 224
rect 198 184 199 224
rect 317 239 318 279
rect 320 239 321 279
rect 1280 11 1320 12
rect 1280 8 1320 9
rect 1380 0 1381 40
rect 1383 0 1384 40
rect 53 -44 93 -43
rect 53 -47 93 -46
rect 153 -55 154 -15
rect 156 -55 157 -15
rect 1280 -40 1320 -39
rect 1280 -43 1320 -42
rect 53 -95 93 -94
rect 53 -98 93 -97
rect 50 -227 51 -187
rect 53 -227 54 -187
rect 77 -227 78 -187
rect 80 -227 81 -187
rect 112 -297 113 -257
rect 115 -297 116 -257
rect 628 -265 629 -225
rect 631 -265 632 -225
rect 655 -265 656 -225
rect 658 -265 659 -225
rect 925 -247 926 -167
rect 928 -247 929 -167
rect 690 -335 691 -295
rect 693 -335 694 -295
rect 925 -347 926 -267
rect 928 -347 929 -267
rect 974 -344 975 -304
rect 977 -344 978 -304
rect 2231 -752 2232 -672
rect 2234 -752 2235 -672
rect 2725 -735 2726 -655
rect 2728 -735 2729 -655
rect 3560 -666 3600 -665
rect 3560 -669 3600 -668
rect 3660 -677 3661 -637
rect 3663 -677 3664 -637
rect 3560 -717 3600 -716
rect 3560 -720 3600 -719
rect 73 -837 113 -836
rect 73 -840 113 -839
rect 173 -848 174 -808
rect 176 -848 177 -808
rect 2231 -852 2232 -772
rect 2234 -852 2235 -772
rect 73 -888 113 -887
rect 73 -891 113 -890
rect 671 -901 672 -861
rect 674 -901 675 -861
rect 698 -901 699 -861
rect 701 -901 702 -861
rect 1009 -910 1010 -870
rect 1012 -910 1013 -870
rect 1036 -910 1037 -870
rect 1039 -910 1040 -870
rect 1389 -899 1390 -859
rect 1392 -899 1393 -859
rect 1416 -899 1417 -859
rect 1419 -899 1420 -859
rect 2280 -849 2281 -809
rect 2283 -849 2284 -809
rect 2725 -835 2726 -755
rect 2728 -835 2729 -755
rect 2774 -832 2775 -792
rect 2777 -832 2778 -792
rect 70 -1020 71 -980
rect 73 -1020 74 -980
rect 97 -1020 98 -980
rect 100 -1020 101 -980
rect 733 -971 734 -931
rect 736 -971 737 -931
rect 1071 -980 1072 -940
rect 1074 -980 1075 -940
rect 1451 -969 1452 -929
rect 1454 -969 1455 -929
rect 132 -1090 133 -1050
rect 135 -1090 136 -1050
rect 5886 -1761 5926 -1760
rect 5886 -1764 5926 -1763
rect 4014 -1859 4015 -1779
rect 4017 -1859 4018 -1779
rect 58 -1961 98 -1960
rect 58 -1964 98 -1963
rect 158 -1972 159 -1932
rect 161 -1972 162 -1932
rect 805 -1962 806 -1922
rect 808 -1962 809 -1922
rect 832 -1962 833 -1922
rect 835 -1962 836 -1922
rect 1273 -1953 1274 -1913
rect 1276 -1953 1277 -1913
rect 1300 -1953 1301 -1913
rect 1303 -1953 1304 -1913
rect 1675 -1950 1676 -1910
rect 1678 -1950 1679 -1910
rect 1702 -1950 1703 -1910
rect 1705 -1950 1706 -1910
rect 2176 -1915 2177 -1875
rect 2179 -1915 2180 -1875
rect 2203 -1915 2204 -1875
rect 2206 -1915 2207 -1875
rect 2781 -1915 2782 -1875
rect 2784 -1915 2785 -1875
rect 2808 -1915 2809 -1875
rect 2811 -1915 2812 -1875
rect 3386 -1915 3387 -1875
rect 3389 -1915 3390 -1875
rect 3413 -1915 3414 -1875
rect 3416 -1915 3417 -1875
rect 58 -2012 98 -2011
rect 58 -2015 98 -2014
rect 867 -2032 868 -1992
rect 870 -2032 871 -1992
rect 1335 -2023 1336 -1983
rect 1338 -2023 1339 -1983
rect 1737 -2020 1738 -1980
rect 1740 -2020 1741 -1980
rect 2238 -1985 2239 -1945
rect 2241 -1985 2242 -1945
rect 2843 -1985 2844 -1945
rect 2846 -1985 2847 -1945
rect 3448 -1985 3449 -1945
rect 3451 -1985 3452 -1945
rect 4014 -1959 4015 -1879
rect 4017 -1959 4018 -1879
rect 4468 -1888 4469 -1808
rect 4471 -1888 4472 -1808
rect 4933 -1853 4934 -1773
rect 4936 -1853 4937 -1773
rect 5986 -1772 5987 -1732
rect 5989 -1772 5990 -1732
rect 5886 -1812 5926 -1811
rect 5886 -1815 5926 -1814
rect 4063 -1956 4064 -1916
rect 4066 -1956 4067 -1916
rect 4468 -1988 4469 -1908
rect 4471 -1988 4472 -1908
rect 4517 -1985 4518 -1945
rect 4520 -1985 4521 -1945
rect 4933 -1953 4934 -1873
rect 4936 -1953 4937 -1873
rect 4982 -1950 4983 -1910
rect 4985 -1950 4986 -1910
rect 55 -2144 56 -2104
rect 58 -2144 59 -2104
rect 82 -2144 83 -2104
rect 85 -2144 86 -2104
rect 117 -2214 118 -2174
rect 120 -2214 121 -2174
rect 6069 -3216 6070 -3136
rect 6072 -3216 6073 -3136
rect 6500 -3210 6501 -3130
rect 6503 -3210 6504 -3130
rect 58 -3380 98 -3379
rect 58 -3383 98 -3382
rect 158 -3391 159 -3351
rect 161 -3391 162 -3351
rect 896 -3388 897 -3348
rect 899 -3388 900 -3348
rect 923 -3388 924 -3348
rect 926 -3388 927 -3348
rect 1234 -3397 1235 -3357
rect 1237 -3397 1238 -3357
rect 1261 -3397 1262 -3357
rect 1264 -3397 1265 -3357
rect 1614 -3386 1615 -3346
rect 1617 -3386 1618 -3346
rect 1641 -3386 1642 -3346
rect 1644 -3386 1645 -3346
rect 2723 -3357 2724 -3317
rect 2726 -3357 2727 -3317
rect 2750 -3357 2751 -3317
rect 2753 -3357 2754 -3317
rect 58 -3431 98 -3430
rect 58 -3434 98 -3433
rect 958 -3458 959 -3418
rect 961 -3458 962 -3418
rect 55 -3563 56 -3523
rect 58 -3563 59 -3523
rect 82 -3563 83 -3523
rect 85 -3563 86 -3523
rect 3061 -3366 3062 -3326
rect 3064 -3366 3065 -3326
rect 3088 -3366 3089 -3326
rect 3091 -3366 3092 -3326
rect 3441 -3355 3442 -3315
rect 3444 -3355 3445 -3315
rect 3468 -3355 3469 -3315
rect 3471 -3355 3472 -3315
rect 4216 -3340 4217 -3300
rect 4219 -3340 4220 -3300
rect 4243 -3340 4244 -3300
rect 4246 -3340 4247 -3300
rect 1296 -3467 1297 -3427
rect 1299 -3467 1300 -3427
rect 1676 -3456 1677 -3416
rect 1679 -3456 1680 -3416
rect 2785 -3427 2786 -3387
rect 2788 -3427 2789 -3387
rect 3123 -3436 3124 -3396
rect 3126 -3436 3127 -3396
rect 4538 -3354 4539 -3314
rect 4541 -3354 4542 -3314
rect 4565 -3354 4566 -3314
rect 4568 -3354 4569 -3314
rect 3503 -3425 3504 -3385
rect 3506 -3425 3507 -3385
rect 4278 -3410 4279 -3370
rect 4281 -3410 4282 -3370
rect 4876 -3363 4877 -3323
rect 4879 -3363 4880 -3323
rect 4903 -3363 4904 -3323
rect 4906 -3363 4907 -3323
rect 5256 -3352 5257 -3312
rect 5259 -3352 5260 -3312
rect 5283 -3352 5284 -3312
rect 5286 -3352 5287 -3312
rect 6069 -3316 6070 -3236
rect 6072 -3316 6073 -3236
rect 6118 -3313 6119 -3273
rect 6121 -3313 6122 -3273
rect 6500 -3310 6501 -3230
rect 6503 -3310 6504 -3230
rect 4600 -3424 4601 -3384
rect 4603 -3424 4604 -3384
rect 6954 -3239 6955 -3159
rect 6957 -3239 6958 -3159
rect 7419 -3204 7420 -3124
rect 7422 -3204 7423 -3124
rect 8560 -3176 8600 -3175
rect 8560 -3179 8600 -3178
rect 8660 -3187 8661 -3147
rect 8663 -3187 8664 -3147
rect 6549 -3307 6550 -3267
rect 6552 -3307 6553 -3267
rect 6954 -3339 6955 -3259
rect 6957 -3339 6958 -3259
rect 7003 -3336 7004 -3296
rect 7006 -3336 7007 -3296
rect 7419 -3304 7420 -3224
rect 7422 -3304 7423 -3224
rect 8560 -3227 8600 -3226
rect 8560 -3230 8600 -3229
rect 7468 -3301 7469 -3261
rect 7471 -3301 7472 -3261
rect 4938 -3433 4939 -3393
rect 4941 -3433 4942 -3393
rect 5318 -3422 5319 -3382
rect 5321 -3422 5322 -3382
rect 117 -3633 118 -3593
rect 120 -3633 121 -3593
<< ndcontact >>
rect -795 546 -775 550
rect -795 538 -775 542
rect -697 531 -693 551
rect -689 531 -685 551
rect -795 495 -775 499
rect -697 498 -693 518
rect -689 498 -685 518
rect -661 496 -657 516
rect -653 496 -649 516
rect -795 487 -775 491
rect -745 288 -741 328
rect -737 288 -733 328
rect -148 306 -128 310
rect -148 298 -128 302
rect -50 291 -46 311
rect -42 291 -38 311
rect -745 223 -741 263
rect -737 223 -733 263
rect -702 254 -698 274
rect -694 254 -690 274
rect -148 255 -128 259
rect -50 258 -46 278
rect -42 258 -38 278
rect -14 256 -10 276
rect -6 256 -2 276
rect -148 247 -128 251
rect 77 240 81 260
rect 85 240 89 260
rect 270 235 274 275
rect 278 235 282 275
rect 270 170 274 210
rect 278 170 282 210
rect 313 201 317 221
rect 321 201 325 221
rect 127 136 131 156
rect 135 136 139 156
rect 160 136 164 156
rect 168 136 172 156
rect 191 146 195 166
rect 199 146 203 166
rect 1242 12 1262 16
rect 1242 4 1262 8
rect 1340 -3 1344 17
rect 1348 -3 1352 17
rect 15 -43 35 -39
rect 15 -51 35 -47
rect 113 -58 117 -38
rect 121 -58 125 -38
rect 1242 -39 1262 -35
rect 1340 -36 1344 -16
rect 1348 -36 1352 -16
rect 1376 -38 1380 -18
rect 1384 -38 1388 -18
rect 1242 -47 1262 -43
rect 15 -94 35 -90
rect 113 -91 117 -71
rect 121 -91 125 -71
rect 149 -93 153 -73
rect 157 -93 161 -73
rect 15 -102 35 -98
rect 65 -301 69 -261
rect 73 -301 77 -261
rect 65 -366 69 -326
rect 73 -366 77 -326
rect 108 -335 112 -315
rect 116 -335 120 -315
rect 643 -339 647 -299
rect 651 -339 655 -299
rect 643 -404 647 -364
rect 651 -404 655 -364
rect 686 -373 690 -353
rect 694 -373 698 -353
rect 906 -392 910 -372
rect 914 -392 918 -372
rect 939 -392 943 -372
rect 947 -392 951 -372
rect 970 -382 974 -362
rect 978 -382 982 -362
rect 3522 -665 3542 -661
rect 3522 -673 3542 -669
rect 3620 -680 3624 -660
rect 3628 -680 3632 -660
rect 3522 -716 3542 -712
rect 3620 -713 3624 -693
rect 3628 -713 3632 -693
rect 3656 -715 3660 -695
rect 3664 -715 3668 -695
rect 3522 -724 3542 -720
rect 35 -836 55 -832
rect 35 -844 55 -840
rect 133 -851 137 -831
rect 141 -851 145 -831
rect 35 -887 55 -883
rect 133 -884 137 -864
rect 141 -884 145 -864
rect 169 -886 173 -866
rect 177 -886 181 -866
rect 35 -895 55 -891
rect 2212 -897 2216 -877
rect 2220 -897 2224 -877
rect 2245 -897 2249 -877
rect 2253 -897 2257 -877
rect 2276 -887 2280 -867
rect 2284 -887 2288 -867
rect 2706 -880 2710 -860
rect 2714 -880 2718 -860
rect 2739 -880 2743 -860
rect 2747 -880 2751 -860
rect 2770 -870 2774 -850
rect 2778 -870 2782 -850
rect 686 -975 690 -935
rect 694 -975 698 -935
rect 1024 -984 1028 -944
rect 1032 -984 1036 -944
rect 85 -1094 89 -1054
rect 93 -1094 97 -1054
rect 686 -1040 690 -1000
rect 694 -1040 698 -1000
rect 729 -1009 733 -989
rect 737 -1009 741 -989
rect 1404 -973 1408 -933
rect 1412 -973 1416 -933
rect 1024 -1049 1028 -1009
rect 1032 -1049 1036 -1009
rect 1067 -1018 1071 -998
rect 1075 -1018 1079 -998
rect 1404 -1038 1408 -998
rect 1412 -1038 1416 -998
rect 1447 -1007 1451 -987
rect 1455 -1007 1459 -987
rect 85 -1159 89 -1119
rect 93 -1159 97 -1119
rect 128 -1128 132 -1108
rect 136 -1128 140 -1108
rect 5848 -1760 5868 -1756
rect 5848 -1768 5868 -1764
rect 20 -1960 40 -1956
rect 20 -1968 40 -1964
rect 118 -1975 122 -1955
rect 126 -1975 130 -1955
rect 20 -2011 40 -2007
rect 118 -2008 122 -1988
rect 126 -2008 130 -1988
rect 154 -2010 158 -1990
rect 162 -2010 166 -1990
rect 20 -2019 40 -2015
rect 820 -2036 824 -1996
rect 828 -2036 832 -1996
rect 1288 -2027 1292 -1987
rect 1296 -2027 1300 -1987
rect 1690 -2024 1694 -1984
rect 1698 -2024 1702 -1984
rect 2191 -1989 2195 -1949
rect 2199 -1989 2203 -1949
rect 2796 -1989 2800 -1949
rect 2804 -1989 2808 -1949
rect 820 -2101 824 -2061
rect 828 -2101 832 -2061
rect 863 -2070 867 -2050
rect 871 -2070 875 -2050
rect 1288 -2092 1292 -2052
rect 1296 -2092 1300 -2052
rect 1331 -2061 1335 -2041
rect 1339 -2061 1343 -2041
rect 1690 -2089 1694 -2049
rect 1698 -2089 1702 -2049
rect 1733 -2058 1737 -2038
rect 1741 -2058 1745 -2038
rect 2191 -2054 2195 -2014
rect 2199 -2054 2203 -2014
rect 2234 -2023 2238 -2003
rect 2242 -2023 2246 -2003
rect 3401 -1989 3405 -1949
rect 3409 -1989 3413 -1949
rect 2796 -2054 2800 -2014
rect 2804 -2054 2808 -2014
rect 2839 -2023 2843 -2003
rect 2847 -2023 2851 -2003
rect 5946 -1775 5950 -1755
rect 5954 -1775 5958 -1755
rect 5848 -1811 5868 -1807
rect 5946 -1808 5950 -1788
rect 5954 -1808 5958 -1788
rect 5982 -1810 5986 -1790
rect 5990 -1810 5994 -1790
rect 5848 -1819 5868 -1815
rect 3401 -2054 3405 -2014
rect 3409 -2054 3413 -2014
rect 3444 -2023 3448 -2003
rect 3452 -2023 3456 -2003
rect 3995 -2004 3999 -1984
rect 4003 -2004 4007 -1984
rect 4028 -2004 4032 -1984
rect 4036 -2004 4040 -1984
rect 4059 -1994 4063 -1974
rect 4067 -1994 4071 -1974
rect 4914 -1998 4918 -1978
rect 4922 -1998 4926 -1978
rect 4947 -1998 4951 -1978
rect 4955 -1998 4959 -1978
rect 4978 -1988 4982 -1968
rect 4986 -1988 4990 -1968
rect 4449 -2033 4453 -2013
rect 4457 -2033 4461 -2013
rect 4482 -2033 4486 -2013
rect 4490 -2033 4494 -2013
rect 4513 -2023 4517 -2003
rect 4521 -2023 4525 -2003
rect 70 -2218 74 -2178
rect 78 -2218 82 -2178
rect 70 -2283 74 -2243
rect 78 -2283 82 -2243
rect 113 -2252 117 -2232
rect 121 -2252 125 -2232
rect 20 -3379 40 -3375
rect 20 -3387 40 -3383
rect 118 -3394 122 -3374
rect 126 -3394 130 -3374
rect 20 -3430 40 -3426
rect 118 -3427 122 -3407
rect 126 -3427 130 -3407
rect 154 -3429 158 -3409
rect 162 -3429 166 -3409
rect 20 -3438 40 -3434
rect 911 -3462 915 -3422
rect 919 -3462 923 -3422
rect 1249 -3471 1253 -3431
rect 1257 -3471 1261 -3431
rect 911 -3527 915 -3487
rect 919 -3527 923 -3487
rect 954 -3496 958 -3476
rect 962 -3496 966 -3476
rect 1629 -3460 1633 -3420
rect 1637 -3460 1641 -3420
rect 2738 -3431 2742 -3391
rect 2746 -3431 2750 -3391
rect 3076 -3440 3080 -3400
rect 3084 -3440 3088 -3400
rect 1249 -3536 1253 -3496
rect 1257 -3536 1261 -3496
rect 1292 -3505 1296 -3485
rect 1300 -3505 1304 -3485
rect 1629 -3525 1633 -3485
rect 1637 -3525 1641 -3485
rect 1672 -3494 1676 -3474
rect 1680 -3494 1684 -3474
rect 2738 -3496 2742 -3456
rect 2746 -3496 2750 -3456
rect 2781 -3465 2785 -3445
rect 2789 -3465 2793 -3445
rect 3456 -3429 3460 -3389
rect 3464 -3429 3468 -3389
rect 4231 -3414 4235 -3374
rect 4239 -3414 4243 -3374
rect 4553 -3428 4557 -3388
rect 4561 -3428 4565 -3388
rect 3076 -3505 3080 -3465
rect 3084 -3505 3088 -3465
rect 3119 -3474 3123 -3454
rect 3127 -3474 3131 -3454
rect 3456 -3494 3460 -3454
rect 3464 -3494 3468 -3454
rect 3499 -3463 3503 -3443
rect 3507 -3463 3511 -3443
rect 4231 -3479 4235 -3439
rect 4239 -3479 4243 -3439
rect 4274 -3448 4278 -3428
rect 4282 -3448 4286 -3428
rect 4891 -3437 4895 -3397
rect 4899 -3437 4903 -3397
rect 4553 -3493 4557 -3453
rect 4561 -3493 4565 -3453
rect 4596 -3462 4600 -3442
rect 4604 -3462 4608 -3442
rect 6050 -3361 6054 -3341
rect 6058 -3361 6062 -3341
rect 6083 -3361 6087 -3341
rect 6091 -3361 6095 -3341
rect 6114 -3351 6118 -3331
rect 6122 -3351 6126 -3331
rect 8522 -3175 8542 -3171
rect 8522 -3183 8542 -3179
rect 8620 -3190 8624 -3170
rect 8628 -3190 8632 -3170
rect 6481 -3355 6485 -3335
rect 6489 -3355 6493 -3335
rect 6514 -3355 6518 -3335
rect 6522 -3355 6526 -3335
rect 6545 -3345 6549 -3325
rect 6553 -3345 6557 -3325
rect 8522 -3226 8542 -3222
rect 8620 -3223 8624 -3203
rect 8628 -3223 8632 -3203
rect 8656 -3225 8660 -3205
rect 8664 -3225 8668 -3205
rect 8522 -3234 8542 -3230
rect 7400 -3349 7404 -3329
rect 7408 -3349 7412 -3329
rect 7433 -3349 7437 -3329
rect 7441 -3349 7445 -3329
rect 7464 -3339 7468 -3319
rect 7472 -3339 7476 -3319
rect 5271 -3426 5275 -3386
rect 5279 -3426 5283 -3386
rect 6935 -3384 6939 -3364
rect 6943 -3384 6947 -3364
rect 6968 -3384 6972 -3364
rect 6976 -3384 6980 -3364
rect 6999 -3374 7003 -3354
rect 7007 -3374 7011 -3354
rect 4891 -3502 4895 -3462
rect 4899 -3502 4903 -3462
rect 4934 -3471 4938 -3451
rect 4942 -3471 4946 -3451
rect 5271 -3491 5275 -3451
rect 5279 -3491 5283 -3451
rect 5314 -3460 5318 -3440
rect 5322 -3460 5326 -3440
rect 70 -3637 74 -3597
rect 78 -3637 82 -3597
rect 70 -3702 74 -3662
rect 78 -3702 82 -3662
rect 113 -3671 117 -3651
rect 121 -3671 125 -3651
<< pdcontact >>
rect -757 546 -717 550
rect -757 538 -717 542
rect -661 534 -657 574
rect -653 534 -649 574
rect -757 495 -717 499
rect -757 487 -717 491
rect -764 362 -760 402
rect -756 362 -752 402
rect -737 362 -733 402
rect -729 362 -725 402
rect -702 292 -698 332
rect -694 292 -690 332
rect -110 306 -70 310
rect -110 298 -70 302
rect -14 294 -10 334
rect -6 294 -2 334
rect -110 255 -70 259
rect 77 278 81 318
rect 85 278 89 318
rect 142 281 146 361
rect 150 281 154 361
rect 251 309 255 349
rect 259 309 263 349
rect 278 309 282 349
rect 286 309 290 349
rect -110 247 -70 251
rect 142 181 146 261
rect 150 181 154 261
rect 191 184 195 224
rect 199 184 203 224
rect 313 239 317 279
rect 321 239 325 279
rect 1280 12 1320 16
rect 1280 4 1320 8
rect 1376 0 1380 40
rect 1384 0 1388 40
rect 53 -43 93 -39
rect 53 -51 93 -47
rect 149 -55 153 -15
rect 157 -55 161 -15
rect 1280 -39 1320 -35
rect 1280 -47 1320 -43
rect 53 -94 93 -90
rect 53 -102 93 -98
rect 46 -227 50 -187
rect 54 -227 58 -187
rect 73 -227 77 -187
rect 81 -227 85 -187
rect 108 -297 112 -257
rect 116 -297 120 -257
rect 624 -265 628 -225
rect 632 -265 636 -225
rect 651 -265 655 -225
rect 659 -265 663 -225
rect 921 -247 925 -167
rect 929 -247 933 -167
rect 686 -335 690 -295
rect 694 -335 698 -295
rect 921 -347 925 -267
rect 929 -347 933 -267
rect 970 -344 974 -304
rect 978 -344 982 -304
rect 2227 -752 2231 -672
rect 2235 -752 2239 -672
rect 2721 -735 2725 -655
rect 2729 -735 2733 -655
rect 3560 -665 3600 -661
rect 3560 -673 3600 -669
rect 3656 -677 3660 -637
rect 3664 -677 3668 -637
rect 3560 -716 3600 -712
rect 3560 -724 3600 -720
rect 73 -836 113 -832
rect 73 -844 113 -840
rect 169 -848 173 -808
rect 177 -848 181 -808
rect 73 -887 113 -883
rect 2227 -852 2231 -772
rect 2235 -852 2239 -772
rect 73 -895 113 -891
rect 667 -901 671 -861
rect 675 -901 679 -861
rect 694 -901 698 -861
rect 702 -901 706 -861
rect 1005 -910 1009 -870
rect 1013 -910 1017 -870
rect 1032 -910 1036 -870
rect 1040 -910 1044 -870
rect 1385 -899 1389 -859
rect 1393 -899 1397 -859
rect 1412 -899 1416 -859
rect 1420 -899 1424 -859
rect 2276 -849 2280 -809
rect 2284 -849 2288 -809
rect 2721 -835 2725 -755
rect 2729 -835 2733 -755
rect 2770 -832 2774 -792
rect 2778 -832 2782 -792
rect 66 -1020 70 -980
rect 74 -1020 78 -980
rect 93 -1020 97 -980
rect 101 -1020 105 -980
rect 729 -971 733 -931
rect 737 -971 741 -931
rect 1067 -980 1071 -940
rect 1075 -980 1079 -940
rect 1447 -969 1451 -929
rect 1455 -969 1459 -929
rect 128 -1090 132 -1050
rect 136 -1090 140 -1050
rect 5886 -1760 5926 -1756
rect 5886 -1768 5926 -1764
rect 4010 -1859 4014 -1779
rect 4018 -1859 4022 -1779
rect 58 -1960 98 -1956
rect 58 -1968 98 -1964
rect 154 -1972 158 -1932
rect 162 -1972 166 -1932
rect 801 -1962 805 -1922
rect 809 -1962 813 -1922
rect 828 -1962 832 -1922
rect 836 -1962 840 -1922
rect 1269 -1953 1273 -1913
rect 1277 -1953 1281 -1913
rect 1296 -1953 1300 -1913
rect 1304 -1953 1308 -1913
rect 1671 -1950 1675 -1910
rect 1679 -1950 1683 -1910
rect 1698 -1950 1702 -1910
rect 1706 -1950 1710 -1910
rect 2172 -1915 2176 -1875
rect 2180 -1915 2184 -1875
rect 2199 -1915 2203 -1875
rect 2207 -1915 2211 -1875
rect 2777 -1915 2781 -1875
rect 2785 -1915 2789 -1875
rect 2804 -1915 2808 -1875
rect 2812 -1915 2816 -1875
rect 3382 -1915 3386 -1875
rect 3390 -1915 3394 -1875
rect 3409 -1915 3413 -1875
rect 3417 -1915 3421 -1875
rect 58 -2011 98 -2007
rect 58 -2019 98 -2015
rect 863 -2032 867 -1992
rect 871 -2032 875 -1992
rect 1331 -2023 1335 -1983
rect 1339 -2023 1343 -1983
rect 1733 -2020 1737 -1980
rect 1741 -2020 1745 -1980
rect 2234 -1985 2238 -1945
rect 2242 -1985 2246 -1945
rect 2839 -1985 2843 -1945
rect 2847 -1985 2851 -1945
rect 3444 -1985 3448 -1945
rect 3452 -1985 3456 -1945
rect 4010 -1959 4014 -1879
rect 4018 -1959 4022 -1879
rect 4464 -1888 4468 -1808
rect 4472 -1888 4476 -1808
rect 4929 -1853 4933 -1773
rect 4937 -1853 4941 -1773
rect 5982 -1772 5986 -1732
rect 5990 -1772 5994 -1732
rect 5886 -1811 5926 -1807
rect 5886 -1819 5926 -1815
rect 4059 -1956 4063 -1916
rect 4067 -1956 4071 -1916
rect 4464 -1988 4468 -1908
rect 4472 -1988 4476 -1908
rect 4513 -1985 4517 -1945
rect 4521 -1985 4525 -1945
rect 4929 -1953 4933 -1873
rect 4937 -1953 4941 -1873
rect 4978 -1950 4982 -1910
rect 4986 -1950 4990 -1910
rect 51 -2144 55 -2104
rect 59 -2144 63 -2104
rect 78 -2144 82 -2104
rect 86 -2144 90 -2104
rect 113 -2214 117 -2174
rect 121 -2214 125 -2174
rect 6065 -3216 6069 -3136
rect 6073 -3216 6077 -3136
rect 6496 -3210 6500 -3130
rect 6504 -3210 6508 -3130
rect 58 -3379 98 -3375
rect 58 -3387 98 -3383
rect 154 -3391 158 -3351
rect 162 -3391 166 -3351
rect 892 -3388 896 -3348
rect 900 -3388 904 -3348
rect 919 -3388 923 -3348
rect 927 -3388 931 -3348
rect 58 -3430 98 -3426
rect 1230 -3397 1234 -3357
rect 1238 -3397 1242 -3357
rect 1257 -3397 1261 -3357
rect 1265 -3397 1269 -3357
rect 1610 -3386 1614 -3346
rect 1618 -3386 1622 -3346
rect 1637 -3386 1641 -3346
rect 1645 -3386 1649 -3346
rect 2719 -3357 2723 -3317
rect 2727 -3357 2731 -3317
rect 2746 -3357 2750 -3317
rect 2754 -3357 2758 -3317
rect 58 -3438 98 -3434
rect 954 -3458 958 -3418
rect 962 -3458 966 -3418
rect 51 -3563 55 -3523
rect 59 -3563 63 -3523
rect 78 -3563 82 -3523
rect 86 -3563 90 -3523
rect 3057 -3366 3061 -3326
rect 3065 -3366 3069 -3326
rect 3084 -3366 3088 -3326
rect 3092 -3366 3096 -3326
rect 3437 -3355 3441 -3315
rect 3445 -3355 3449 -3315
rect 3464 -3355 3468 -3315
rect 3472 -3355 3476 -3315
rect 4212 -3340 4216 -3300
rect 4220 -3340 4224 -3300
rect 4239 -3340 4243 -3300
rect 4247 -3340 4251 -3300
rect 1292 -3467 1296 -3427
rect 1300 -3467 1304 -3427
rect 1672 -3456 1676 -3416
rect 1680 -3456 1684 -3416
rect 2781 -3427 2785 -3387
rect 2789 -3427 2793 -3387
rect 3119 -3436 3123 -3396
rect 3127 -3436 3131 -3396
rect 4534 -3354 4538 -3314
rect 4542 -3354 4546 -3314
rect 4561 -3354 4565 -3314
rect 4569 -3354 4573 -3314
rect 3499 -3425 3503 -3385
rect 3507 -3425 3511 -3385
rect 4274 -3410 4278 -3370
rect 4282 -3410 4286 -3370
rect 4872 -3363 4876 -3323
rect 4880 -3363 4884 -3323
rect 4899 -3363 4903 -3323
rect 4907 -3363 4911 -3323
rect 5252 -3352 5256 -3312
rect 5260 -3352 5264 -3312
rect 5279 -3352 5283 -3312
rect 5287 -3352 5291 -3312
rect 6065 -3316 6069 -3236
rect 6073 -3316 6077 -3236
rect 6114 -3313 6118 -3273
rect 6122 -3313 6126 -3273
rect 6496 -3310 6500 -3230
rect 6504 -3310 6508 -3230
rect 4596 -3424 4600 -3384
rect 4604 -3424 4608 -3384
rect 6950 -3239 6954 -3159
rect 6958 -3239 6962 -3159
rect 7415 -3204 7419 -3124
rect 7423 -3204 7427 -3124
rect 8560 -3175 8600 -3171
rect 8560 -3183 8600 -3179
rect 8656 -3187 8660 -3147
rect 8664 -3187 8668 -3147
rect 6545 -3307 6549 -3267
rect 6553 -3307 6557 -3267
rect 6950 -3339 6954 -3259
rect 6958 -3339 6962 -3259
rect 6999 -3336 7003 -3296
rect 7007 -3336 7011 -3296
rect 7415 -3304 7419 -3224
rect 7423 -3304 7427 -3224
rect 8560 -3226 8600 -3222
rect 8560 -3234 8600 -3230
rect 7464 -3301 7468 -3261
rect 7472 -3301 7476 -3261
rect 4934 -3433 4938 -3393
rect 4942 -3433 4946 -3393
rect 5314 -3422 5318 -3382
rect 5322 -3422 5326 -3382
rect 113 -3633 117 -3593
rect 121 -3633 125 -3593
<< psubstratepcontact >>
rect -806 553 -802 557
rect -806 532 -802 536
rect -806 502 -802 506
rect -806 481 -802 485
rect -668 485 -664 489
rect -647 485 -643 489
rect -159 313 -155 317
rect -159 292 -155 296
rect -159 262 -155 266
rect -709 243 -705 247
rect -688 243 -684 247
rect -159 241 -155 245
rect -21 245 -17 249
rect 0 245 4 249
rect 70 229 74 233
rect 91 229 95 233
rect -752 212 -748 216
rect -731 212 -727 216
rect 306 190 310 194
rect 327 190 331 194
rect 263 159 267 163
rect 284 159 288 163
rect 184 135 188 139
rect 205 135 209 139
rect 120 125 124 129
rect 141 125 145 129
rect 153 125 157 129
rect 174 125 178 129
rect 1231 19 1235 23
rect 1231 -2 1235 2
rect 4 -36 8 -32
rect 4 -57 8 -53
rect 1231 -32 1235 -28
rect 1231 -53 1235 -49
rect 1369 -49 1373 -45
rect 1390 -49 1394 -45
rect 4 -87 8 -83
rect 4 -108 8 -104
rect 142 -104 146 -100
rect 163 -104 167 -100
rect 101 -346 105 -342
rect 122 -346 126 -342
rect 58 -377 62 -373
rect 79 -377 83 -373
rect 679 -384 683 -380
rect 700 -384 704 -380
rect 963 -393 967 -389
rect 984 -393 988 -389
rect 899 -403 903 -399
rect 920 -403 924 -399
rect 932 -403 936 -399
rect 953 -403 957 -399
rect 636 -415 640 -411
rect 657 -415 661 -411
rect 3511 -658 3515 -654
rect 3511 -679 3515 -675
rect 3511 -709 3515 -705
rect 3511 -730 3515 -726
rect 3649 -726 3653 -722
rect 3670 -726 3674 -722
rect 24 -829 28 -825
rect 24 -850 28 -846
rect 24 -880 28 -876
rect 24 -901 28 -897
rect 162 -897 166 -893
rect 183 -897 187 -893
rect 2763 -881 2767 -877
rect 2784 -881 2788 -877
rect 2699 -891 2703 -887
rect 2720 -891 2724 -887
rect 2732 -891 2736 -887
rect 2753 -891 2757 -887
rect 2269 -898 2273 -894
rect 2290 -898 2294 -894
rect 2205 -908 2209 -904
rect 2226 -908 2230 -904
rect 2238 -908 2242 -904
rect 2259 -908 2263 -904
rect 722 -1020 726 -1016
rect 743 -1020 747 -1016
rect 679 -1051 683 -1047
rect 700 -1051 704 -1047
rect 1060 -1029 1064 -1025
rect 1081 -1029 1085 -1025
rect 1440 -1018 1444 -1014
rect 1461 -1018 1465 -1014
rect 1397 -1049 1401 -1045
rect 1418 -1049 1422 -1045
rect 1017 -1060 1021 -1056
rect 1038 -1060 1042 -1056
rect 121 -1139 125 -1135
rect 142 -1139 146 -1135
rect 78 -1170 82 -1166
rect 99 -1170 103 -1166
rect 5837 -1753 5841 -1749
rect 9 -1953 13 -1949
rect 9 -1974 13 -1970
rect 9 -2004 13 -2000
rect 9 -2025 13 -2021
rect 147 -2021 151 -2017
rect 168 -2021 172 -2017
rect 856 -2081 860 -2077
rect 877 -2081 881 -2077
rect 1324 -2072 1328 -2068
rect 1345 -2072 1349 -2068
rect 2227 -2034 2231 -2030
rect 2248 -2034 2252 -2030
rect 5837 -1774 5841 -1770
rect 5837 -1804 5841 -1800
rect 5837 -1825 5841 -1821
rect 5975 -1821 5979 -1817
rect 5996 -1821 6000 -1817
rect 2832 -2034 2836 -2030
rect 2853 -2034 2857 -2030
rect 4052 -2005 4056 -2001
rect 4073 -2005 4077 -2001
rect 3988 -2015 3992 -2011
rect 4009 -2015 4013 -2011
rect 4021 -2015 4025 -2011
rect 4042 -2015 4046 -2011
rect 4971 -1999 4975 -1995
rect 4992 -1999 4996 -1995
rect 3437 -2034 3441 -2030
rect 3458 -2034 3462 -2030
rect 4907 -2009 4911 -2005
rect 4928 -2009 4932 -2005
rect 4940 -2009 4944 -2005
rect 4961 -2009 4965 -2005
rect 4506 -2034 4510 -2030
rect 4527 -2034 4531 -2030
rect 4442 -2044 4446 -2040
rect 4463 -2044 4467 -2040
rect 4475 -2044 4479 -2040
rect 4496 -2044 4500 -2040
rect 2184 -2065 2188 -2061
rect 2205 -2065 2209 -2061
rect 2789 -2065 2793 -2061
rect 2810 -2065 2814 -2061
rect 3394 -2065 3398 -2061
rect 3415 -2065 3419 -2061
rect 1726 -2069 1730 -2065
rect 1747 -2069 1751 -2065
rect 1281 -2103 1285 -2099
rect 1302 -2103 1306 -2099
rect 1683 -2100 1687 -2096
rect 1704 -2100 1708 -2096
rect 813 -2112 817 -2108
rect 834 -2112 838 -2108
rect 106 -2263 110 -2259
rect 127 -2263 131 -2259
rect 63 -2294 67 -2290
rect 84 -2294 88 -2290
rect 9 -3372 13 -3368
rect 9 -3393 13 -3389
rect 9 -3423 13 -3419
rect 9 -3444 13 -3440
rect 147 -3440 151 -3436
rect 168 -3440 172 -3436
rect 947 -3507 951 -3503
rect 968 -3507 972 -3503
rect 904 -3538 908 -3534
rect 925 -3538 929 -3534
rect 1285 -3516 1289 -3512
rect 1306 -3516 1310 -3512
rect 2774 -3476 2778 -3472
rect 2795 -3476 2799 -3472
rect 1665 -3505 1669 -3501
rect 1686 -3505 1690 -3501
rect 2731 -3507 2735 -3503
rect 2752 -3507 2756 -3503
rect 3112 -3485 3116 -3481
rect 3133 -3485 3137 -3481
rect 3492 -3474 3496 -3470
rect 3513 -3474 3517 -3470
rect 4267 -3459 4271 -3455
rect 4288 -3459 4292 -3455
rect 4224 -3490 4228 -3486
rect 4245 -3490 4249 -3486
rect 8511 -3168 8515 -3164
rect 8511 -3189 8515 -3185
rect 6538 -3356 6542 -3352
rect 6559 -3356 6563 -3352
rect 6107 -3362 6111 -3358
rect 6128 -3362 6132 -3358
rect 6474 -3366 6478 -3362
rect 6495 -3366 6499 -3362
rect 6507 -3366 6511 -3362
rect 6528 -3366 6532 -3362
rect 8511 -3219 8515 -3215
rect 8511 -3240 8515 -3236
rect 8649 -3236 8653 -3232
rect 8670 -3236 8674 -3232
rect 7457 -3350 7461 -3346
rect 7478 -3350 7482 -3346
rect 6043 -3372 6047 -3368
rect 6064 -3372 6068 -3368
rect 6076 -3372 6080 -3368
rect 6097 -3372 6101 -3368
rect 7393 -3360 7397 -3356
rect 7414 -3360 7418 -3356
rect 7426 -3360 7430 -3356
rect 7447 -3360 7451 -3356
rect 6992 -3385 6996 -3381
rect 7013 -3385 7017 -3381
rect 6928 -3395 6932 -3391
rect 6949 -3395 6953 -3391
rect 6961 -3395 6965 -3391
rect 6982 -3395 6986 -3391
rect 4589 -3473 4593 -3469
rect 4610 -3473 4614 -3469
rect 3449 -3505 3453 -3501
rect 3470 -3505 3474 -3501
rect 4546 -3504 4550 -3500
rect 4567 -3504 4571 -3500
rect 4927 -3482 4931 -3478
rect 4948 -3482 4952 -3478
rect 5307 -3471 5311 -3467
rect 5328 -3471 5332 -3467
rect 5264 -3502 5268 -3498
rect 5285 -3502 5289 -3498
rect 3069 -3516 3073 -3512
rect 3090 -3516 3094 -3512
rect 4884 -3513 4888 -3509
rect 4905 -3513 4909 -3509
rect 1622 -3536 1626 -3532
rect 1643 -3536 1647 -3532
rect 1242 -3547 1246 -3543
rect 1263 -3547 1267 -3543
rect 106 -3682 110 -3678
rect 127 -3682 131 -3678
rect 63 -3713 67 -3709
rect 84 -3713 88 -3709
<< nsubstratencontact >>
rect -666 581 -662 585
rect -649 581 -645 585
rect -710 551 -706 555
rect -710 534 -706 538
rect -710 500 -706 504
rect -710 483 -706 487
rect -769 409 -765 413
rect -752 409 -748 413
rect -742 409 -738 413
rect -725 409 -721 413
rect 137 368 141 372
rect 154 368 158 372
rect -707 339 -703 343
rect -690 339 -686 343
rect -19 341 -15 345
rect -2 341 2 345
rect -63 311 -59 315
rect -63 294 -59 298
rect 72 325 76 329
rect 89 325 93 329
rect -63 260 -59 264
rect 246 356 250 360
rect 263 356 267 360
rect 273 356 277 360
rect 290 356 294 360
rect -63 243 -59 247
rect 186 231 190 235
rect 203 231 207 235
rect 308 286 312 290
rect 325 286 329 290
rect 1371 47 1375 51
rect 1388 47 1392 51
rect 1327 17 1331 21
rect 1327 0 1331 4
rect 144 -8 148 -4
rect 161 -8 165 -4
rect 100 -38 104 -34
rect 100 -55 104 -51
rect 1327 -34 1331 -30
rect 1327 -51 1331 -47
rect 100 -89 104 -85
rect 100 -106 104 -102
rect 916 -160 920 -156
rect 933 -160 937 -156
rect 41 -180 45 -176
rect 58 -180 62 -176
rect 68 -180 72 -176
rect 85 -180 89 -176
rect 619 -218 623 -214
rect 636 -218 640 -214
rect 646 -218 650 -214
rect 663 -218 667 -214
rect 103 -250 107 -246
rect 120 -250 124 -246
rect 681 -288 685 -284
rect 698 -288 702 -284
rect 965 -297 969 -293
rect 982 -297 986 -293
rect 3651 -630 3655 -626
rect 3668 -630 3672 -626
rect 2716 -648 2720 -644
rect 2733 -648 2737 -644
rect 2222 -665 2226 -661
rect 2239 -665 2243 -661
rect 3607 -660 3611 -656
rect 3607 -677 3611 -673
rect 3607 -711 3611 -707
rect 3607 -728 3611 -724
rect 164 -801 168 -797
rect 181 -801 185 -797
rect 120 -831 124 -827
rect 120 -848 124 -844
rect 120 -882 124 -878
rect 662 -854 666 -850
rect 679 -854 683 -850
rect 689 -854 693 -850
rect 706 -854 710 -850
rect 1380 -852 1384 -848
rect 1397 -852 1401 -848
rect 1407 -852 1411 -848
rect 1424 -852 1428 -848
rect 120 -899 124 -895
rect 1000 -863 1004 -859
rect 1017 -863 1021 -859
rect 1027 -863 1031 -859
rect 1044 -863 1048 -859
rect 2271 -802 2275 -798
rect 2288 -802 2292 -798
rect 2765 -785 2769 -781
rect 2782 -785 2786 -781
rect 61 -973 65 -969
rect 78 -973 82 -969
rect 88 -973 92 -969
rect 105 -973 109 -969
rect 724 -924 728 -920
rect 741 -924 745 -920
rect 123 -1043 127 -1039
rect 140 -1043 144 -1039
rect 1062 -933 1066 -929
rect 1079 -933 1083 -929
rect 1442 -922 1446 -918
rect 1459 -922 1463 -918
rect 5977 -1725 5981 -1721
rect 5994 -1725 5998 -1721
rect 5933 -1755 5937 -1751
rect 4924 -1766 4928 -1762
rect 4941 -1766 4945 -1762
rect 4005 -1772 4009 -1768
rect 4022 -1772 4026 -1768
rect 4459 -1801 4463 -1797
rect 4476 -1801 4480 -1797
rect 2167 -1868 2171 -1864
rect 2184 -1868 2188 -1864
rect 2194 -1868 2198 -1864
rect 2211 -1868 2215 -1864
rect 2772 -1868 2776 -1864
rect 2789 -1868 2793 -1864
rect 2799 -1868 2803 -1864
rect 2816 -1868 2820 -1864
rect 3377 -1868 3381 -1864
rect 3394 -1868 3398 -1864
rect 3404 -1868 3408 -1864
rect 3421 -1868 3425 -1864
rect 1264 -1906 1268 -1902
rect 1281 -1906 1285 -1902
rect 1291 -1906 1295 -1902
rect 1308 -1906 1312 -1902
rect 1666 -1903 1670 -1899
rect 1683 -1903 1687 -1899
rect 1693 -1903 1697 -1899
rect 1710 -1903 1714 -1899
rect 796 -1915 800 -1911
rect 813 -1915 817 -1911
rect 823 -1915 827 -1911
rect 840 -1915 844 -1911
rect 149 -1925 153 -1921
rect 166 -1925 170 -1921
rect 105 -1955 109 -1951
rect 105 -1972 109 -1968
rect 105 -2006 109 -2002
rect 105 -2023 109 -2019
rect 858 -1985 862 -1981
rect 875 -1985 879 -1981
rect 1326 -1976 1330 -1972
rect 1343 -1976 1347 -1972
rect 1728 -1973 1732 -1969
rect 1745 -1973 1749 -1969
rect 2229 -1938 2233 -1934
rect 2246 -1938 2250 -1934
rect 46 -2097 50 -2093
rect 63 -2097 67 -2093
rect 73 -2097 77 -2093
rect 90 -2097 94 -2093
rect 2834 -1938 2838 -1934
rect 2851 -1938 2855 -1934
rect 3439 -1938 3443 -1934
rect 3456 -1938 3460 -1934
rect 5933 -1772 5937 -1768
rect 5933 -1806 5937 -1802
rect 5933 -1823 5937 -1819
rect 4054 -1909 4058 -1905
rect 4071 -1909 4075 -1905
rect 4508 -1938 4512 -1934
rect 4525 -1938 4529 -1934
rect 4973 -1903 4977 -1899
rect 4990 -1903 4994 -1899
rect 108 -2167 112 -2163
rect 125 -2167 129 -2163
rect 7410 -3117 7414 -3113
rect 7427 -3117 7431 -3113
rect 6491 -3123 6495 -3119
rect 6508 -3123 6512 -3119
rect 6060 -3129 6064 -3125
rect 6077 -3129 6081 -3125
rect 6945 -3152 6949 -3148
rect 6962 -3152 6966 -3148
rect 4207 -3293 4211 -3289
rect 4224 -3293 4228 -3289
rect 4234 -3293 4238 -3289
rect 4251 -3293 4255 -3289
rect 2714 -3310 2718 -3306
rect 2731 -3310 2735 -3306
rect 2741 -3310 2745 -3306
rect 2758 -3310 2762 -3306
rect 3432 -3308 3436 -3304
rect 3449 -3308 3453 -3304
rect 3459 -3308 3463 -3304
rect 3476 -3308 3480 -3304
rect 149 -3344 153 -3340
rect 166 -3344 170 -3340
rect 887 -3341 891 -3337
rect 904 -3341 908 -3337
rect 914 -3341 918 -3337
rect 931 -3341 935 -3337
rect 1605 -3339 1609 -3335
rect 1622 -3339 1626 -3335
rect 1632 -3339 1636 -3335
rect 1649 -3339 1653 -3335
rect 105 -3374 109 -3370
rect 105 -3391 109 -3387
rect 1225 -3350 1229 -3346
rect 1242 -3350 1246 -3346
rect 1252 -3350 1256 -3346
rect 1269 -3350 1273 -3346
rect 105 -3425 109 -3421
rect 3052 -3319 3056 -3315
rect 3069 -3319 3073 -3315
rect 3079 -3319 3083 -3315
rect 3096 -3319 3100 -3315
rect 105 -3442 109 -3438
rect 949 -3411 953 -3407
rect 966 -3411 970 -3407
rect 46 -3516 50 -3512
rect 63 -3516 67 -3512
rect 73 -3516 77 -3512
rect 90 -3516 94 -3512
rect 4529 -3307 4533 -3303
rect 4546 -3307 4550 -3303
rect 4556 -3307 4560 -3303
rect 4573 -3307 4577 -3303
rect 5247 -3305 5251 -3301
rect 5264 -3305 5268 -3301
rect 5274 -3305 5278 -3301
rect 5291 -3305 5295 -3301
rect 1287 -3420 1291 -3416
rect 1304 -3420 1308 -3416
rect 1667 -3409 1671 -3405
rect 1684 -3409 1688 -3405
rect 2776 -3380 2780 -3376
rect 2793 -3380 2797 -3376
rect 3114 -3389 3118 -3385
rect 3131 -3389 3135 -3385
rect 4867 -3316 4871 -3312
rect 4884 -3316 4888 -3312
rect 4894 -3316 4898 -3312
rect 4911 -3316 4915 -3312
rect 3494 -3378 3498 -3374
rect 3511 -3378 3515 -3374
rect 4269 -3363 4273 -3359
rect 4286 -3363 4290 -3359
rect 6109 -3266 6113 -3262
rect 6126 -3266 6130 -3262
rect 4591 -3377 4595 -3373
rect 4608 -3377 4612 -3373
rect 8651 -3140 8655 -3136
rect 8668 -3140 8672 -3136
rect 8607 -3170 8611 -3166
rect 8607 -3187 8611 -3183
rect 6540 -3260 6544 -3256
rect 6557 -3260 6561 -3256
rect 6994 -3289 6998 -3285
rect 7011 -3289 7015 -3285
rect 8607 -3221 8611 -3217
rect 8607 -3238 8611 -3234
rect 7459 -3254 7463 -3250
rect 7476 -3254 7480 -3250
rect 4929 -3386 4933 -3382
rect 4946 -3386 4950 -3382
rect 5309 -3375 5313 -3371
rect 5326 -3375 5330 -3371
rect 108 -3586 112 -3582
rect 125 -3586 129 -3582
<< polysilicon >>
rect -772 573 -690 575
rect -656 574 -654 577
rect -692 551 -690 573
rect -798 543 -795 545
rect -775 543 -757 545
rect -717 543 -714 545
rect -692 528 -690 531
rect -772 521 -690 523
rect -692 518 -690 521
rect -656 516 -654 534
rect -692 495 -690 498
rect -798 492 -795 494
rect -775 492 -757 494
rect -717 492 -714 494
rect -656 493 -654 496
rect -759 402 -757 405
rect -732 402 -730 405
rect -759 334 -757 362
rect -732 350 -730 362
rect 147 361 149 364
rect -732 348 -722 350
rect -759 332 -738 334
rect -740 328 -738 332
rect -740 284 -738 288
rect -724 271 -722 348
rect -697 332 -695 335
rect -125 333 -43 335
rect -9 334 -7 337
rect -45 311 -43 333
rect -151 303 -148 305
rect -128 303 -110 305
rect -70 303 -67 305
rect -697 274 -695 292
rect 82 318 84 321
rect -45 288 -43 291
rect -125 281 -43 283
rect -45 278 -43 281
rect -740 269 -722 271
rect -740 263 -738 269
rect -9 276 -7 294
rect 256 349 258 352
rect 283 349 285 352
rect -45 255 -43 258
rect 82 260 84 278
rect 147 275 149 281
rect 256 281 258 309
rect 283 297 285 309
rect 283 295 293 297
rect 256 279 277 281
rect 275 275 277 279
rect 147 273 167 275
rect 147 261 149 264
rect -697 251 -695 254
rect -151 252 -148 254
rect -128 252 -110 254
rect -70 252 -67 254
rect -9 253 -7 256
rect 82 237 84 240
rect -740 220 -738 223
rect 147 175 149 181
rect 132 173 149 175
rect 132 156 134 173
rect 165 156 167 273
rect 275 231 277 235
rect 196 224 198 227
rect 291 218 293 295
rect 318 279 320 282
rect 318 221 320 239
rect 275 216 293 218
rect 275 210 277 216
rect 196 166 198 184
rect 318 198 320 201
rect 275 167 277 170
rect 196 143 198 146
rect 132 133 134 136
rect 165 133 167 136
rect 1265 39 1347 41
rect 1381 40 1383 43
rect 1345 17 1347 39
rect 1239 9 1242 11
rect 1262 9 1280 11
rect 1320 9 1323 11
rect 1345 -6 1347 -3
rect 38 -16 120 -14
rect 154 -15 156 -12
rect 1265 -13 1347 -11
rect 118 -38 120 -16
rect 12 -46 15 -44
rect 35 -46 53 -44
rect 93 -46 96 -44
rect 1345 -16 1347 -13
rect 1381 -18 1383 0
rect 1345 -39 1347 -36
rect 1239 -42 1242 -40
rect 1262 -42 1280 -40
rect 1320 -42 1323 -40
rect 1381 -41 1383 -38
rect 118 -61 120 -58
rect 38 -68 120 -66
rect 118 -71 120 -68
rect 154 -73 156 -55
rect 118 -94 120 -91
rect 12 -97 15 -95
rect 35 -97 53 -95
rect 93 -97 96 -95
rect 154 -96 156 -93
rect 926 -167 928 -164
rect 51 -187 53 -184
rect 78 -187 80 -184
rect 629 -225 631 -222
rect 656 -225 658 -222
rect 51 -255 53 -227
rect 78 -239 80 -227
rect 78 -241 88 -239
rect 51 -257 72 -255
rect 70 -261 72 -257
rect 70 -305 72 -301
rect 86 -318 88 -241
rect 113 -257 115 -254
rect 926 -253 928 -247
rect 926 -255 946 -253
rect 629 -293 631 -265
rect 656 -277 658 -265
rect 926 -267 928 -264
rect 656 -279 666 -277
rect 629 -295 650 -293
rect 113 -315 115 -297
rect 648 -299 650 -295
rect 70 -320 88 -318
rect 70 -326 72 -320
rect 113 -338 115 -335
rect 648 -343 650 -339
rect 664 -356 666 -279
rect 691 -295 693 -292
rect 691 -353 693 -335
rect 926 -353 928 -347
rect 648 -358 666 -356
rect 648 -364 650 -358
rect 70 -369 72 -366
rect 911 -355 928 -353
rect 911 -372 913 -355
rect 944 -372 946 -255
rect 975 -304 977 -301
rect 975 -362 977 -344
rect 691 -376 693 -373
rect 975 -385 977 -382
rect 911 -395 913 -392
rect 944 -395 946 -392
rect 648 -407 650 -404
rect 3545 -638 3627 -636
rect 3661 -637 3663 -634
rect 2726 -655 2728 -652
rect 2232 -672 2234 -669
rect 3625 -660 3627 -638
rect 3519 -668 3522 -666
rect 3542 -668 3560 -666
rect 3600 -668 3603 -666
rect 3625 -683 3627 -680
rect 3545 -690 3627 -688
rect 3625 -693 3627 -690
rect 3661 -695 3663 -677
rect 3625 -716 3627 -713
rect 3519 -719 3522 -717
rect 3542 -719 3560 -717
rect 3600 -719 3603 -717
rect 3661 -718 3663 -715
rect 2726 -741 2728 -735
rect 2726 -743 2746 -741
rect 2232 -758 2234 -752
rect 2726 -755 2728 -752
rect 2232 -760 2252 -758
rect 2232 -772 2234 -769
rect 58 -809 140 -807
rect 174 -808 176 -805
rect 138 -831 140 -809
rect 32 -839 35 -837
rect 55 -839 73 -837
rect 113 -839 116 -837
rect 138 -854 140 -851
rect 58 -861 140 -859
rect 138 -864 140 -861
rect 174 -866 176 -848
rect 672 -861 674 -858
rect 699 -861 701 -858
rect 1390 -859 1392 -856
rect 1417 -859 1419 -856
rect 2232 -858 2234 -852
rect 138 -887 140 -884
rect 32 -890 35 -888
rect 55 -890 73 -888
rect 113 -890 116 -888
rect 174 -889 176 -886
rect 1010 -870 1012 -867
rect 1037 -870 1039 -867
rect 672 -929 674 -901
rect 699 -913 701 -901
rect 2217 -860 2234 -858
rect 2217 -877 2219 -860
rect 2250 -877 2252 -760
rect 2281 -809 2283 -806
rect 2726 -841 2728 -835
rect 2711 -843 2728 -841
rect 2281 -867 2283 -849
rect 2711 -860 2713 -843
rect 2744 -860 2746 -743
rect 2775 -792 2777 -789
rect 2775 -850 2777 -832
rect 2775 -873 2777 -870
rect 2711 -883 2713 -880
rect 2744 -883 2746 -880
rect 2281 -890 2283 -887
rect 699 -915 709 -913
rect 672 -931 693 -929
rect 691 -935 693 -931
rect 71 -980 73 -977
rect 98 -980 100 -977
rect 691 -979 693 -975
rect 707 -992 709 -915
rect 734 -931 736 -928
rect 1010 -938 1012 -910
rect 1037 -922 1039 -910
rect 1037 -924 1047 -922
rect 1010 -940 1031 -938
rect 1029 -944 1031 -940
rect 734 -989 736 -971
rect 1029 -988 1031 -984
rect 691 -994 709 -992
rect 691 -1000 693 -994
rect 71 -1048 73 -1020
rect 98 -1032 100 -1020
rect 98 -1034 108 -1032
rect 71 -1050 92 -1048
rect 90 -1054 92 -1050
rect 90 -1098 92 -1094
rect 106 -1111 108 -1034
rect 1045 -1001 1047 -924
rect 1390 -927 1392 -899
rect 1417 -911 1419 -899
rect 2217 -900 2219 -897
rect 2250 -900 2252 -897
rect 1417 -913 1427 -911
rect 1390 -929 1411 -927
rect 1409 -933 1411 -929
rect 1072 -940 1074 -937
rect 1409 -977 1411 -973
rect 1072 -998 1074 -980
rect 1425 -990 1427 -913
rect 1452 -929 1454 -926
rect 1452 -987 1454 -969
rect 1409 -992 1427 -990
rect 1409 -998 1411 -992
rect 1029 -1003 1047 -1001
rect 1029 -1009 1031 -1003
rect 734 -1012 736 -1009
rect 691 -1043 693 -1040
rect 133 -1050 135 -1047
rect 1072 -1021 1074 -1018
rect 1452 -1010 1454 -1007
rect 1409 -1041 1411 -1038
rect 1029 -1052 1031 -1049
rect 133 -1108 135 -1090
rect 90 -1113 108 -1111
rect 90 -1119 92 -1113
rect 133 -1131 135 -1128
rect 90 -1162 92 -1159
rect 5871 -1733 5953 -1731
rect 5987 -1732 5989 -1729
rect 5951 -1755 5953 -1733
rect 5845 -1763 5848 -1761
rect 5868 -1763 5886 -1761
rect 5926 -1763 5929 -1761
rect 4934 -1773 4936 -1770
rect 4015 -1779 4017 -1776
rect 4469 -1808 4471 -1805
rect 4015 -1865 4017 -1859
rect 4015 -1867 4035 -1865
rect 2177 -1875 2179 -1872
rect 2204 -1875 2206 -1872
rect 2782 -1875 2784 -1872
rect 2809 -1875 2811 -1872
rect 3387 -1875 3389 -1872
rect 3414 -1875 3416 -1872
rect 1676 -1910 1678 -1907
rect 1703 -1910 1705 -1907
rect 1274 -1913 1276 -1910
rect 1301 -1913 1303 -1910
rect 806 -1922 808 -1919
rect 833 -1922 835 -1919
rect 43 -1933 125 -1931
rect 159 -1932 161 -1929
rect 123 -1955 125 -1933
rect 17 -1963 20 -1961
rect 40 -1963 58 -1961
rect 98 -1963 101 -1961
rect 4015 -1879 4017 -1876
rect 2177 -1943 2179 -1915
rect 2204 -1927 2206 -1915
rect 2204 -1929 2214 -1927
rect 2177 -1945 2198 -1943
rect 2196 -1949 2198 -1945
rect 123 -1978 125 -1975
rect 43 -1985 125 -1983
rect 123 -1988 125 -1985
rect 159 -1990 161 -1972
rect 123 -2011 125 -2008
rect 806 -1990 808 -1962
rect 833 -1974 835 -1962
rect 833 -1976 843 -1974
rect 806 -1992 827 -1990
rect 825 -1996 827 -1992
rect 17 -2014 20 -2012
rect 40 -2014 58 -2012
rect 98 -2014 101 -2012
rect 159 -2013 161 -2010
rect 825 -2040 827 -2036
rect 841 -2053 843 -1976
rect 1274 -1981 1276 -1953
rect 1301 -1965 1303 -1953
rect 1301 -1967 1311 -1965
rect 1274 -1983 1295 -1981
rect 1293 -1987 1295 -1983
rect 868 -1992 870 -1989
rect 1293 -2031 1295 -2027
rect 868 -2050 870 -2032
rect 1309 -2044 1311 -1967
rect 1676 -1978 1678 -1950
rect 1703 -1962 1705 -1950
rect 1703 -1964 1713 -1962
rect 1676 -1980 1697 -1978
rect 1336 -1983 1338 -1980
rect 1695 -1984 1697 -1980
rect 1336 -2041 1338 -2023
rect 1695 -2028 1697 -2024
rect 1711 -2041 1713 -1964
rect 1738 -1980 1740 -1977
rect 2196 -1993 2198 -1989
rect 2212 -2006 2214 -1929
rect 2239 -1945 2241 -1942
rect 2782 -1943 2784 -1915
rect 2809 -1927 2811 -1915
rect 2809 -1929 2819 -1927
rect 2782 -1945 2803 -1943
rect 2801 -1949 2803 -1945
rect 2239 -2003 2241 -1985
rect 2801 -1993 2803 -1989
rect 2196 -2008 2214 -2006
rect 2196 -2014 2198 -2008
rect 1738 -2038 1740 -2020
rect 1293 -2046 1311 -2044
rect 825 -2055 843 -2053
rect 825 -2061 827 -2055
rect 1293 -2052 1295 -2046
rect 868 -2073 870 -2070
rect 1695 -2043 1713 -2041
rect 1695 -2049 1697 -2043
rect 1336 -2064 1338 -2061
rect 2817 -2006 2819 -1929
rect 2844 -1945 2846 -1942
rect 3387 -1943 3389 -1915
rect 3414 -1927 3416 -1915
rect 3414 -1929 3424 -1927
rect 3387 -1945 3408 -1943
rect 3406 -1949 3408 -1945
rect 2844 -2003 2846 -1985
rect 3406 -1993 3408 -1989
rect 2801 -2008 2819 -2006
rect 2801 -2014 2803 -2008
rect 2239 -2026 2241 -2023
rect 3422 -2006 3424 -1929
rect 3449 -1945 3451 -1942
rect 4015 -1965 4017 -1959
rect 4000 -1967 4017 -1965
rect 4000 -1984 4002 -1967
rect 4033 -1984 4035 -1867
rect 5951 -1778 5953 -1775
rect 5871 -1785 5953 -1783
rect 5951 -1788 5953 -1785
rect 5987 -1790 5989 -1772
rect 5951 -1811 5953 -1808
rect 5845 -1814 5848 -1812
rect 5868 -1814 5886 -1812
rect 5926 -1814 5929 -1812
rect 5987 -1813 5989 -1810
rect 4934 -1859 4936 -1853
rect 4934 -1861 4954 -1859
rect 4934 -1873 4936 -1870
rect 4469 -1894 4471 -1888
rect 4469 -1896 4489 -1894
rect 4469 -1908 4471 -1905
rect 4064 -1916 4066 -1913
rect 4064 -1974 4066 -1956
rect 3449 -2003 3451 -1985
rect 3406 -2008 3424 -2006
rect 3406 -2014 3408 -2008
rect 2844 -2026 2846 -2023
rect 4469 -1994 4471 -1988
rect 4064 -1997 4066 -1994
rect 4454 -1996 4471 -1994
rect 4000 -2007 4002 -2004
rect 4033 -2007 4035 -2004
rect 4454 -2013 4456 -1996
rect 4487 -2013 4489 -1896
rect 4518 -1945 4520 -1942
rect 4934 -1959 4936 -1953
rect 4919 -1961 4936 -1959
rect 4919 -1978 4921 -1961
rect 4952 -1978 4954 -1861
rect 4983 -1910 4985 -1907
rect 4983 -1968 4985 -1950
rect 4518 -2003 4520 -1985
rect 4983 -1991 4985 -1988
rect 4919 -2001 4921 -1998
rect 4952 -2001 4954 -1998
rect 3449 -2026 3451 -2023
rect 4518 -2026 4520 -2023
rect 4454 -2036 4456 -2033
rect 4487 -2036 4489 -2033
rect 2196 -2057 2198 -2054
rect 2801 -2057 2803 -2054
rect 3406 -2057 3408 -2054
rect 1738 -2061 1740 -2058
rect 1695 -2092 1697 -2089
rect 1293 -2095 1295 -2092
rect 56 -2104 58 -2101
rect 83 -2104 85 -2101
rect 825 -2104 827 -2101
rect 56 -2172 58 -2144
rect 83 -2156 85 -2144
rect 83 -2158 93 -2156
rect 56 -2174 77 -2172
rect 75 -2178 77 -2174
rect 75 -2222 77 -2218
rect 91 -2235 93 -2158
rect 118 -2174 120 -2171
rect 118 -2232 120 -2214
rect 75 -2237 93 -2235
rect 75 -2243 77 -2237
rect 118 -2255 120 -2252
rect 75 -2286 77 -2283
rect 7420 -3124 7422 -3121
rect 6501 -3130 6503 -3127
rect 6070 -3136 6072 -3133
rect 6955 -3159 6957 -3156
rect 6070 -3222 6072 -3216
rect 6501 -3216 6503 -3210
rect 6501 -3218 6521 -3216
rect 6070 -3224 6090 -3222
rect 6070 -3236 6072 -3233
rect 4217 -3300 4219 -3297
rect 4244 -3300 4246 -3297
rect 2724 -3317 2726 -3314
rect 2751 -3317 2753 -3314
rect 3442 -3315 3444 -3312
rect 3469 -3315 3471 -3312
rect 897 -3348 899 -3345
rect 924 -3348 926 -3345
rect 1615 -3346 1617 -3343
rect 1642 -3346 1644 -3343
rect 43 -3352 125 -3350
rect 159 -3351 161 -3348
rect 123 -3374 125 -3352
rect 17 -3382 20 -3380
rect 40 -3382 58 -3380
rect 98 -3382 101 -3380
rect 1235 -3357 1237 -3354
rect 1262 -3357 1264 -3354
rect 123 -3397 125 -3394
rect 43 -3404 125 -3402
rect 123 -3407 125 -3404
rect 159 -3409 161 -3391
rect 123 -3430 125 -3427
rect 897 -3416 899 -3388
rect 924 -3400 926 -3388
rect 3062 -3326 3064 -3323
rect 3089 -3326 3091 -3323
rect 924 -3402 934 -3400
rect 897 -3418 918 -3416
rect 916 -3422 918 -3418
rect 17 -3433 20 -3431
rect 40 -3433 58 -3431
rect 98 -3433 101 -3431
rect 159 -3432 161 -3429
rect 916 -3466 918 -3462
rect 932 -3479 934 -3402
rect 959 -3418 961 -3415
rect 1235 -3425 1237 -3397
rect 1262 -3409 1264 -3397
rect 1262 -3411 1272 -3409
rect 1235 -3427 1256 -3425
rect 1254 -3431 1256 -3427
rect 959 -3476 961 -3458
rect 1254 -3475 1256 -3471
rect 916 -3481 934 -3479
rect 916 -3487 918 -3481
rect 56 -3523 58 -3520
rect 83 -3523 85 -3520
rect 1270 -3488 1272 -3411
rect 1615 -3414 1617 -3386
rect 1642 -3398 1644 -3386
rect 2724 -3385 2726 -3357
rect 2751 -3369 2753 -3357
rect 4539 -3314 4541 -3311
rect 4566 -3314 4568 -3311
rect 5257 -3312 5259 -3309
rect 5284 -3312 5286 -3309
rect 2751 -3371 2761 -3369
rect 2724 -3387 2745 -3385
rect 2743 -3391 2745 -3387
rect 1642 -3400 1652 -3398
rect 1615 -3416 1636 -3414
rect 1634 -3420 1636 -3416
rect 1297 -3427 1299 -3424
rect 1634 -3464 1636 -3460
rect 1297 -3485 1299 -3467
rect 1650 -3477 1652 -3400
rect 1677 -3416 1679 -3413
rect 2743 -3435 2745 -3431
rect 2759 -3448 2761 -3371
rect 2786 -3387 2788 -3384
rect 3062 -3394 3064 -3366
rect 3089 -3378 3091 -3366
rect 3089 -3380 3099 -3378
rect 3062 -3396 3083 -3394
rect 3081 -3400 3083 -3396
rect 2786 -3445 2788 -3427
rect 3081 -3444 3083 -3440
rect 2743 -3450 2761 -3448
rect 2743 -3456 2745 -3450
rect 1677 -3474 1679 -3456
rect 1634 -3479 1652 -3477
rect 1634 -3485 1636 -3479
rect 1254 -3490 1272 -3488
rect 1254 -3496 1256 -3490
rect 959 -3499 961 -3496
rect 916 -3530 918 -3527
rect 1297 -3508 1299 -3505
rect 1677 -3497 1679 -3494
rect 3097 -3457 3099 -3380
rect 3442 -3383 3444 -3355
rect 3469 -3367 3471 -3355
rect 3469 -3369 3479 -3367
rect 3442 -3385 3463 -3383
rect 3461 -3389 3463 -3385
rect 3124 -3396 3126 -3393
rect 3461 -3433 3463 -3429
rect 3124 -3454 3126 -3436
rect 3477 -3446 3479 -3369
rect 4217 -3368 4219 -3340
rect 4244 -3352 4246 -3340
rect 4244 -3354 4254 -3352
rect 4877 -3323 4879 -3320
rect 4904 -3323 4906 -3320
rect 4217 -3370 4238 -3368
rect 4236 -3374 4238 -3370
rect 3504 -3385 3506 -3382
rect 4236 -3418 4238 -3414
rect 3504 -3443 3506 -3425
rect 4252 -3431 4254 -3354
rect 4279 -3370 4281 -3367
rect 4539 -3382 4541 -3354
rect 4566 -3366 4568 -3354
rect 6070 -3322 6072 -3316
rect 6055 -3324 6072 -3322
rect 6055 -3341 6057 -3324
rect 6088 -3341 6090 -3224
rect 6501 -3230 6503 -3227
rect 6119 -3273 6121 -3270
rect 6119 -3331 6121 -3313
rect 6501 -3316 6503 -3310
rect 6486 -3318 6503 -3316
rect 4566 -3368 4576 -3366
rect 4539 -3384 4560 -3382
rect 4558 -3388 4560 -3384
rect 4279 -3428 4281 -3410
rect 4236 -3433 4254 -3431
rect 4236 -3439 4238 -3433
rect 3461 -3448 3479 -3446
rect 3461 -3454 3463 -3448
rect 3081 -3459 3099 -3457
rect 3081 -3465 3083 -3459
rect 2786 -3468 2788 -3465
rect 2743 -3499 2745 -3496
rect 3124 -3477 3126 -3474
rect 3504 -3466 3506 -3463
rect 4558 -3432 4560 -3428
rect 4574 -3445 4576 -3368
rect 4601 -3384 4603 -3381
rect 4877 -3391 4879 -3363
rect 4904 -3375 4906 -3363
rect 4904 -3377 4914 -3375
rect 4877 -3393 4898 -3391
rect 4896 -3397 4898 -3393
rect 4601 -3442 4603 -3424
rect 4896 -3441 4898 -3437
rect 4279 -3451 4281 -3448
rect 4558 -3447 4576 -3445
rect 4558 -3453 4560 -3447
rect 4236 -3482 4238 -3479
rect 4912 -3454 4914 -3377
rect 5257 -3380 5259 -3352
rect 5284 -3364 5286 -3352
rect 6486 -3335 6488 -3318
rect 6519 -3335 6521 -3218
rect 8545 -3148 8627 -3146
rect 8661 -3147 8663 -3144
rect 8625 -3170 8627 -3148
rect 8519 -3178 8522 -3176
rect 8542 -3178 8560 -3176
rect 8600 -3178 8603 -3176
rect 8625 -3193 8627 -3190
rect 8545 -3200 8627 -3198
rect 8625 -3203 8627 -3200
rect 7420 -3210 7422 -3204
rect 7420 -3212 7440 -3210
rect 7420 -3224 7422 -3221
rect 6955 -3245 6957 -3239
rect 6955 -3247 6975 -3245
rect 6955 -3259 6957 -3256
rect 6550 -3267 6552 -3264
rect 6550 -3325 6552 -3307
rect 6119 -3354 6121 -3351
rect 6955 -3345 6957 -3339
rect 6550 -3348 6552 -3345
rect 6940 -3347 6957 -3345
rect 6486 -3358 6488 -3355
rect 6519 -3358 6521 -3355
rect 6055 -3364 6057 -3361
rect 6088 -3364 6090 -3361
rect 5284 -3366 5294 -3364
rect 6940 -3364 6942 -3347
rect 6973 -3364 6975 -3247
rect 7004 -3296 7006 -3293
rect 7420 -3310 7422 -3304
rect 7405 -3312 7422 -3310
rect 7405 -3329 7407 -3312
rect 7438 -3329 7440 -3212
rect 8661 -3205 8663 -3187
rect 8625 -3226 8627 -3223
rect 8519 -3229 8522 -3227
rect 8542 -3229 8560 -3227
rect 8600 -3229 8603 -3227
rect 8661 -3228 8663 -3225
rect 7469 -3261 7471 -3258
rect 7469 -3319 7471 -3301
rect 7004 -3354 7006 -3336
rect 7469 -3342 7471 -3339
rect 7405 -3352 7407 -3349
rect 7438 -3352 7440 -3349
rect 5257 -3382 5278 -3380
rect 5276 -3386 5278 -3382
rect 4939 -3393 4941 -3390
rect 5276 -3430 5278 -3426
rect 4939 -3451 4941 -3433
rect 5292 -3443 5294 -3366
rect 5319 -3382 5321 -3379
rect 7004 -3377 7006 -3374
rect 6940 -3387 6942 -3384
rect 6973 -3387 6975 -3384
rect 5319 -3440 5321 -3422
rect 5276 -3445 5294 -3443
rect 5276 -3451 5278 -3445
rect 4896 -3456 4914 -3454
rect 4896 -3462 4898 -3456
rect 4601 -3465 4603 -3462
rect 3461 -3497 3463 -3494
rect 4558 -3496 4560 -3493
rect 4939 -3474 4941 -3471
rect 5319 -3463 5321 -3460
rect 5276 -3494 5278 -3491
rect 4896 -3505 4898 -3502
rect 3081 -3508 3083 -3505
rect 1634 -3528 1636 -3525
rect 1254 -3539 1256 -3536
rect 56 -3591 58 -3563
rect 83 -3575 85 -3563
rect 83 -3577 93 -3575
rect 56 -3593 77 -3591
rect 75 -3597 77 -3593
rect 75 -3641 77 -3637
rect 91 -3654 93 -3577
rect 118 -3593 120 -3590
rect 118 -3651 120 -3633
rect 75 -3656 93 -3654
rect 75 -3662 77 -3656
rect 118 -3674 120 -3671
rect 75 -3705 77 -3702
<< polycontact >>
rect -772 568 -767 573
rect -772 545 -767 550
rect -772 523 -767 528
rect -661 519 -656 524
rect -772 494 -767 499
rect -764 332 -759 337
rect -125 328 -120 333
rect -125 305 -120 310
rect -702 277 -697 282
rect -125 283 -120 288
rect -14 279 -9 284
rect -745 266 -740 271
rect -125 254 -120 259
rect 77 263 82 268
rect 142 273 147 278
rect 251 279 256 284
rect 127 170 132 175
rect 313 224 318 229
rect 270 213 275 218
rect 191 169 196 174
rect 1265 34 1270 39
rect 1265 11 1270 16
rect 1265 -11 1270 -6
rect 38 -21 43 -16
rect 38 -44 43 -39
rect 1376 -15 1381 -10
rect 1265 -40 1270 -35
rect 38 -66 43 -61
rect 149 -70 154 -65
rect 38 -95 43 -90
rect 46 -257 51 -252
rect 921 -255 926 -250
rect 624 -295 629 -290
rect 108 -312 113 -307
rect 65 -323 70 -318
rect 686 -350 691 -345
rect 643 -361 648 -356
rect 906 -358 911 -353
rect 970 -359 975 -354
rect 3545 -643 3550 -638
rect 3545 -666 3550 -661
rect 3545 -688 3550 -683
rect 3656 -692 3661 -687
rect 3545 -717 3550 -712
rect 2721 -743 2726 -738
rect 2227 -760 2232 -755
rect 58 -814 63 -809
rect 58 -837 63 -832
rect 58 -859 63 -854
rect 169 -863 174 -858
rect 58 -888 63 -883
rect 667 -931 672 -926
rect 2212 -863 2217 -858
rect 2706 -846 2711 -841
rect 2276 -864 2281 -859
rect 2770 -847 2775 -842
rect 1005 -940 1010 -935
rect 729 -986 734 -981
rect 686 -997 691 -992
rect 66 -1050 71 -1045
rect 1385 -929 1390 -924
rect 1067 -995 1072 -990
rect 1447 -984 1452 -979
rect 1404 -995 1409 -990
rect 1024 -1006 1029 -1001
rect 128 -1105 133 -1100
rect 85 -1116 90 -1111
rect 5871 -1738 5876 -1733
rect 5871 -1761 5876 -1756
rect 4010 -1867 4015 -1862
rect 43 -1938 48 -1933
rect 43 -1961 48 -1956
rect 2172 -1945 2177 -1940
rect 43 -1983 48 -1978
rect 154 -1987 159 -1982
rect 43 -2012 48 -2007
rect 801 -1992 806 -1987
rect 1269 -1983 1274 -1978
rect 863 -2047 868 -2042
rect 1671 -1980 1676 -1975
rect 1331 -2038 1336 -2033
rect 2777 -1945 2782 -1940
rect 2234 -2000 2239 -1995
rect 2191 -2011 2196 -2006
rect 1733 -2035 1738 -2030
rect 1288 -2049 1293 -2044
rect 820 -2058 825 -2053
rect 1690 -2046 1695 -2041
rect 3382 -1945 3387 -1940
rect 2839 -2000 2844 -1995
rect 2796 -2011 2801 -2006
rect 3995 -1970 4000 -1965
rect 5871 -1783 5876 -1778
rect 5982 -1787 5987 -1782
rect 5871 -1812 5876 -1807
rect 4929 -1861 4934 -1856
rect 4464 -1896 4469 -1891
rect 4059 -1971 4064 -1966
rect 3444 -2000 3449 -1995
rect 3401 -2011 3406 -2006
rect 4449 -1999 4454 -1994
rect 4914 -1964 4919 -1959
rect 4978 -1965 4983 -1960
rect 4513 -2000 4518 -1995
rect 51 -2174 56 -2169
rect 113 -2229 118 -2224
rect 70 -2240 75 -2235
rect 6065 -3224 6070 -3219
rect 6496 -3218 6501 -3213
rect 43 -3357 48 -3352
rect 43 -3380 48 -3375
rect 43 -3402 48 -3397
rect 154 -3406 159 -3401
rect 43 -3431 48 -3426
rect 892 -3418 897 -3413
rect 1230 -3427 1235 -3422
rect 954 -3473 959 -3468
rect 911 -3484 916 -3479
rect 1610 -3416 1615 -3411
rect 2719 -3387 2724 -3382
rect 1292 -3482 1297 -3477
rect 3057 -3396 3062 -3391
rect 2781 -3442 2786 -3437
rect 2738 -3453 2743 -3448
rect 1672 -3471 1677 -3466
rect 1629 -3482 1634 -3477
rect 1249 -3493 1254 -3488
rect 3437 -3385 3442 -3380
rect 3119 -3451 3124 -3446
rect 4212 -3370 4217 -3365
rect 3499 -3440 3504 -3435
rect 4534 -3384 4539 -3379
rect 6050 -3327 6055 -3322
rect 6114 -3328 6119 -3323
rect 6481 -3321 6486 -3316
rect 4274 -3425 4279 -3420
rect 4231 -3436 4236 -3431
rect 3456 -3451 3461 -3446
rect 3076 -3462 3081 -3457
rect 4872 -3393 4877 -3388
rect 4596 -3439 4601 -3434
rect 4553 -3450 4558 -3445
rect 5252 -3382 5257 -3377
rect 8545 -3153 8550 -3148
rect 8545 -3176 8550 -3171
rect 8545 -3198 8550 -3193
rect 8656 -3202 8661 -3197
rect 7415 -3212 7420 -3207
rect 6950 -3247 6955 -3242
rect 6545 -3322 6550 -3317
rect 6935 -3350 6940 -3345
rect 7400 -3315 7405 -3310
rect 8545 -3227 8550 -3222
rect 7464 -3316 7469 -3311
rect 6999 -3351 7004 -3346
rect 4934 -3448 4939 -3443
rect 5314 -3437 5319 -3432
rect 5271 -3448 5276 -3443
rect 4891 -3459 4896 -3454
rect 51 -3593 56 -3588
rect 113 -3648 118 -3643
rect 70 -3659 75 -3654
<< metal1 >>
rect -669 585 -642 588
rect -669 581 -666 585
rect -662 581 -649 585
rect -645 581 -642 585
rect -669 579 -642 581
rect -661 574 -657 579
rect -772 566 -767 568
rect -904 561 -767 566
rect -867 271 -858 561
rect -807 557 -801 558
rect -807 553 -806 557
rect -802 553 -801 557
rect -807 550 -801 553
rect -772 550 -767 561
rect -712 555 -703 558
rect -712 551 -710 555
rect -706 551 -703 555
rect -689 551 -676 554
rect -712 550 -703 551
rect -807 546 -795 550
rect -807 536 -801 546
rect -717 546 -703 550
rect -775 538 -757 542
rect -712 538 -703 546
rect -807 532 -806 536
rect -802 532 -801 536
rect -807 531 -801 532
rect -772 528 -767 538
rect -712 534 -710 538
rect -706 534 -703 538
rect -712 531 -703 534
rect -697 528 -693 531
rect -743 524 -693 528
rect -743 519 -739 524
rect -833 514 -739 519
rect -689 518 -685 531
rect -682 524 -676 551
rect -653 524 -649 534
rect -682 519 -661 524
rect -653 519 -642 524
rect -842 337 -833 514
rect -807 506 -801 507
rect -807 502 -806 506
rect -802 502 -801 506
rect -807 499 -801 502
rect -772 499 -767 514
rect -712 504 -703 507
rect -712 500 -710 504
rect -706 500 -703 504
rect -712 499 -703 500
rect -807 495 -795 499
rect -807 485 -801 495
rect -717 495 -703 499
rect -775 487 -757 491
rect -712 487 -703 495
rect -807 481 -806 485
rect -802 481 -801 485
rect -807 480 -801 481
rect -772 467 -767 487
rect -712 483 -710 487
rect -706 483 -703 487
rect -712 480 -703 483
rect -653 516 -649 519
rect -697 467 -693 498
rect -661 490 -657 496
rect -669 489 -642 490
rect -669 485 -668 489
rect -664 485 -647 489
rect -643 485 -642 489
rect -669 484 -642 485
rect -772 464 -693 467
rect -772 413 -718 416
rect -772 409 -769 413
rect -765 409 -752 413
rect -748 409 -742 413
rect -738 409 -725 413
rect -721 409 -718 413
rect -772 407 -718 409
rect -764 402 -760 407
rect -737 402 -733 407
rect 134 372 161 375
rect 134 368 137 372
rect 141 368 154 372
rect 158 368 161 372
rect 134 366 161 368
rect -756 342 -752 362
rect -729 342 -725 362
rect 142 361 146 366
rect -710 343 -683 346
rect -756 338 -715 342
rect -842 332 -764 337
rect -842 331 -833 332
rect -737 328 -733 338
rect -745 282 -741 288
rect -720 282 -715 338
rect -710 339 -707 343
rect -703 339 -690 343
rect -686 339 -683 343
rect -22 345 5 348
rect -22 341 -19 345
rect -15 341 -2 345
rect 2 341 5 345
rect -22 339 5 341
rect -710 337 -683 339
rect -702 332 -698 337
rect -14 334 -10 339
rect -125 326 -120 328
rect -160 321 -120 326
rect -694 282 -690 292
rect -160 317 -154 318
rect -160 313 -159 317
rect -155 313 -154 317
rect -160 310 -154 313
rect -125 310 -120 321
rect -65 315 -56 318
rect -65 311 -63 315
rect -59 311 -56 315
rect -42 311 -29 314
rect -65 310 -56 311
rect -160 306 -148 310
rect -160 296 -154 306
rect -70 306 -56 310
rect -128 298 -110 302
rect -65 298 -56 306
rect -160 292 -159 296
rect -155 292 -154 296
rect -160 291 -154 292
rect -125 288 -120 298
rect -65 294 -63 298
rect -59 294 -56 298
rect -65 291 -56 294
rect -50 288 -46 291
rect -96 284 -46 288
rect -745 278 -731 282
rect -737 277 -731 278
rect -720 277 -702 282
rect -694 277 -681 282
rect -96 279 -92 284
rect -867 266 -745 271
rect -737 263 -733 277
rect -694 274 -690 277
rect -160 274 -92 279
rect -42 278 -38 291
rect -35 284 -29 311
rect 69 329 96 332
rect 69 325 72 329
rect 76 325 89 329
rect 93 325 96 329
rect 69 323 96 325
rect -6 284 -2 294
rect 77 318 81 323
rect -35 279 -14 284
rect -6 279 5 284
rect -160 266 -154 267
rect -160 262 -159 266
rect -155 262 -154 266
rect -160 259 -154 262
rect -125 259 -120 274
rect -65 264 -56 267
rect -65 260 -63 264
rect -59 260 -56 264
rect -65 259 -56 260
rect -160 255 -148 259
rect -702 248 -698 254
rect -710 247 -683 248
rect -710 243 -709 247
rect -705 243 -688 247
rect -684 243 -683 247
rect -710 242 -683 243
rect -160 245 -154 255
rect -70 255 -56 259
rect -128 247 -110 251
rect -65 247 -56 255
rect -160 241 -159 245
rect -155 241 -154 245
rect -160 240 -154 241
rect -125 227 -120 247
rect -65 243 -63 247
rect -59 243 -56 247
rect -65 240 -56 243
rect -6 276 -2 279
rect 243 360 297 363
rect 243 356 246 360
rect 250 356 263 360
rect 267 356 273 360
rect 277 356 290 360
rect 294 356 297 360
rect 243 354 297 356
rect 251 349 255 354
rect 278 349 282 354
rect 259 289 263 309
rect 286 289 290 309
rect 305 290 332 293
rect 259 285 300 289
rect -50 227 -46 258
rect 85 268 89 278
rect 125 273 142 278
rect 150 269 154 281
rect 244 279 251 284
rect 278 275 282 285
rect 69 263 77 268
rect 85 263 98 268
rect 142 265 154 269
rect 85 260 89 263
rect -14 250 -10 256
rect -22 249 5 250
rect -22 245 -21 249
rect -17 245 0 249
rect 4 245 5 249
rect -22 244 5 245
rect 142 261 146 265
rect 77 234 81 240
rect 69 233 96 234
rect 69 229 70 233
rect 74 229 91 233
rect 95 229 96 233
rect 69 228 96 229
rect -125 224 -46 227
rect -745 217 -741 223
rect -753 216 -726 217
rect -753 212 -752 216
rect -748 212 -731 216
rect -727 212 -726 216
rect -753 211 -726 212
rect 183 235 210 238
rect 183 231 186 235
rect 190 231 203 235
rect 207 231 210 235
rect 183 229 210 231
rect 270 229 274 235
rect 295 229 300 285
rect 305 286 308 290
rect 312 286 325 290
rect 329 286 332 290
rect 305 284 332 286
rect 313 279 317 284
rect 321 229 325 239
rect 191 224 195 229
rect 270 225 284 229
rect 278 224 284 225
rect 295 224 313 229
rect 321 224 334 229
rect 244 213 270 218
rect 278 210 282 224
rect 321 221 325 224
rect 118 170 127 175
rect 150 174 154 181
rect 199 174 203 184
rect 150 169 191 174
rect 199 169 210 174
rect 313 195 317 201
rect 305 194 332 195
rect 305 190 306 194
rect 310 190 327 194
rect 331 190 332 194
rect 305 189 332 190
rect 150 166 154 169
rect 199 166 203 169
rect 135 162 172 166
rect 135 156 139 162
rect 168 156 172 162
rect 270 164 274 170
rect 262 163 289 164
rect 262 159 263 163
rect 267 159 284 163
rect 288 159 289 163
rect 262 158 289 159
rect 191 140 195 146
rect 183 139 210 140
rect 127 130 131 136
rect 160 130 164 136
rect 183 135 184 139
rect 188 135 205 139
rect 209 135 210 139
rect 183 134 210 135
rect 119 129 146 130
rect 119 125 120 129
rect 124 125 141 129
rect 145 125 146 129
rect 119 124 146 125
rect 152 129 179 130
rect 152 125 153 129
rect 157 125 174 129
rect 178 125 179 129
rect 152 124 179 125
rect 1368 51 1395 54
rect 1368 47 1371 51
rect 1375 47 1388 51
rect 1392 47 1395 51
rect 1368 45 1395 47
rect 1376 40 1380 45
rect 1265 32 1270 34
rect 1230 27 1270 32
rect 1230 23 1236 24
rect 1230 19 1231 23
rect 1235 19 1236 23
rect 1230 16 1236 19
rect 1265 16 1270 27
rect 1325 21 1334 24
rect 1325 17 1327 21
rect 1331 17 1334 21
rect 1348 17 1361 20
rect 1325 16 1334 17
rect 1230 12 1242 16
rect 1230 2 1236 12
rect 1320 12 1334 16
rect 1262 4 1280 8
rect 1325 4 1334 12
rect 141 -4 168 -1
rect 1230 -2 1231 2
rect 1235 -2 1236 2
rect 1230 -3 1236 -2
rect 141 -8 144 -4
rect 148 -8 161 -4
rect 165 -8 168 -4
rect 141 -10 168 -8
rect 1265 -6 1270 4
rect 1325 0 1327 4
rect 1331 0 1334 4
rect 1325 -3 1334 0
rect 1340 -6 1344 -3
rect 149 -15 153 -10
rect 1294 -10 1344 -6
rect 1294 -15 1298 -10
rect 38 -23 43 -21
rect -94 -28 43 -23
rect -57 -318 -48 -28
rect 3 -32 9 -31
rect 3 -36 4 -32
rect 8 -36 9 -32
rect 3 -39 9 -36
rect 38 -39 43 -28
rect 98 -34 107 -31
rect 98 -38 100 -34
rect 104 -38 107 -34
rect 121 -38 134 -35
rect 98 -39 107 -38
rect 3 -43 15 -39
rect 3 -53 9 -43
rect 93 -43 107 -39
rect 35 -51 53 -47
rect 98 -51 107 -43
rect 3 -57 4 -53
rect 8 -57 9 -53
rect 3 -58 9 -57
rect 38 -61 43 -51
rect 98 -55 100 -51
rect 104 -55 107 -51
rect 98 -58 107 -55
rect 113 -61 117 -58
rect 67 -65 117 -61
rect 67 -70 71 -65
rect -23 -75 71 -70
rect 121 -71 125 -58
rect 128 -65 134 -38
rect 1230 -20 1298 -15
rect 1348 -16 1352 -3
rect 1355 -10 1361 17
rect 1384 -10 1388 0
rect 1355 -15 1376 -10
rect 1384 -15 1395 -10
rect 1230 -28 1236 -27
rect 1230 -32 1231 -28
rect 1235 -32 1236 -28
rect 1230 -35 1236 -32
rect 1265 -35 1270 -20
rect 1325 -30 1334 -27
rect 1325 -34 1327 -30
rect 1331 -34 1334 -30
rect 1325 -35 1334 -34
rect 1230 -39 1242 -35
rect 1230 -49 1236 -39
rect 1320 -39 1334 -35
rect 1262 -47 1280 -43
rect 1325 -47 1334 -39
rect 1230 -53 1231 -49
rect 1235 -53 1236 -49
rect 1230 -54 1236 -53
rect 157 -65 161 -55
rect 128 -70 149 -65
rect 157 -70 168 -65
rect 1265 -67 1270 -47
rect 1325 -51 1327 -47
rect 1331 -51 1334 -47
rect 1325 -54 1334 -51
rect 1384 -18 1388 -15
rect 1340 -67 1344 -36
rect 1376 -44 1380 -38
rect 1368 -45 1395 -44
rect 1368 -49 1369 -45
rect 1373 -49 1390 -45
rect 1394 -49 1395 -45
rect 1368 -50 1395 -49
rect 1265 -70 1344 -67
rect -32 -252 -23 -75
rect 3 -83 9 -82
rect 3 -87 4 -83
rect 8 -87 9 -83
rect 3 -90 9 -87
rect 38 -90 43 -75
rect 98 -85 107 -82
rect 98 -89 100 -85
rect 104 -89 107 -85
rect 98 -90 107 -89
rect 3 -94 15 -90
rect 3 -104 9 -94
rect 93 -94 107 -90
rect 35 -102 53 -98
rect 98 -102 107 -94
rect 3 -108 4 -104
rect 8 -108 9 -104
rect 3 -109 9 -108
rect 38 -122 43 -102
rect 98 -106 100 -102
rect 104 -106 107 -102
rect 98 -109 107 -106
rect 157 -73 161 -70
rect 113 -122 117 -91
rect 149 -99 153 -93
rect 141 -100 168 -99
rect 141 -104 142 -100
rect 146 -104 163 -100
rect 167 -104 168 -100
rect 141 -105 168 -104
rect 38 -125 117 -122
rect 913 -156 940 -153
rect 913 -160 916 -156
rect 920 -160 933 -156
rect 937 -160 940 -156
rect 913 -162 940 -160
rect 921 -167 925 -162
rect 38 -176 92 -173
rect 38 -180 41 -176
rect 45 -180 58 -176
rect 62 -180 68 -176
rect 72 -180 85 -176
rect 89 -180 92 -176
rect 38 -182 92 -180
rect 46 -187 50 -182
rect 73 -187 77 -182
rect 616 -214 670 -211
rect 616 -218 619 -214
rect 623 -218 636 -214
rect 640 -218 646 -214
rect 650 -218 663 -214
rect 667 -218 670 -214
rect 616 -220 670 -218
rect 54 -247 58 -227
rect 81 -247 85 -227
rect 624 -225 628 -220
rect 651 -225 655 -220
rect 100 -246 127 -243
rect 54 -251 95 -247
rect -32 -257 46 -252
rect -32 -258 -23 -257
rect 73 -261 77 -251
rect 65 -307 69 -301
rect 90 -307 95 -251
rect 100 -250 103 -246
rect 107 -250 120 -246
rect 124 -250 127 -246
rect 100 -252 127 -250
rect 108 -257 112 -252
rect 904 -255 921 -250
rect 929 -259 933 -247
rect 632 -285 636 -265
rect 659 -285 663 -265
rect 921 -263 933 -259
rect 921 -267 925 -263
rect 678 -284 705 -281
rect 632 -289 673 -285
rect 617 -295 624 -290
rect 116 -307 120 -297
rect 651 -299 655 -289
rect 65 -311 79 -307
rect 73 -312 79 -311
rect 90 -312 108 -307
rect 116 -312 129 -307
rect -57 -323 65 -318
rect 73 -326 77 -312
rect 116 -315 120 -312
rect 108 -341 112 -335
rect 100 -342 127 -341
rect 100 -346 101 -342
rect 105 -346 122 -342
rect 126 -346 127 -342
rect 100 -347 127 -346
rect 643 -345 647 -339
rect 668 -345 673 -289
rect 678 -288 681 -284
rect 685 -288 698 -284
rect 702 -288 705 -284
rect 678 -290 705 -288
rect 686 -295 690 -290
rect 694 -345 698 -335
rect 643 -349 657 -345
rect 651 -350 657 -349
rect 668 -350 686 -345
rect 694 -350 707 -345
rect 962 -293 989 -290
rect 962 -297 965 -293
rect 969 -297 982 -293
rect 986 -297 989 -293
rect 962 -299 989 -297
rect 970 -304 974 -299
rect 617 -361 643 -356
rect 651 -364 655 -350
rect 694 -353 698 -350
rect 65 -372 69 -366
rect 57 -373 84 -372
rect 57 -377 58 -373
rect 62 -377 79 -373
rect 83 -377 84 -373
rect 57 -378 84 -377
rect 897 -358 906 -353
rect 929 -354 933 -347
rect 978 -354 982 -344
rect 929 -359 970 -354
rect 978 -359 989 -354
rect 929 -362 933 -359
rect 978 -362 982 -359
rect 914 -366 951 -362
rect 914 -372 918 -366
rect 947 -372 951 -366
rect 686 -379 690 -373
rect 678 -380 705 -379
rect 678 -384 679 -380
rect 683 -384 700 -380
rect 704 -384 705 -380
rect 678 -385 705 -384
rect 970 -388 974 -382
rect 962 -389 989 -388
rect 906 -398 910 -392
rect 939 -398 943 -392
rect 962 -393 963 -389
rect 967 -393 984 -389
rect 988 -393 989 -389
rect 962 -394 989 -393
rect 898 -399 925 -398
rect 898 -403 899 -399
rect 903 -403 920 -399
rect 924 -403 925 -399
rect 898 -404 925 -403
rect 931 -399 958 -398
rect 931 -403 932 -399
rect 936 -403 953 -399
rect 957 -403 958 -399
rect 931 -404 958 -403
rect 643 -410 647 -404
rect 635 -411 662 -410
rect 635 -415 636 -411
rect 640 -415 657 -411
rect 661 -415 662 -411
rect 635 -416 662 -415
rect 3648 -626 3675 -623
rect 3648 -630 3651 -626
rect 3655 -630 3668 -626
rect 3672 -630 3675 -626
rect 3648 -632 3675 -630
rect 3656 -637 3660 -632
rect 2713 -644 2740 -641
rect 2713 -648 2716 -644
rect 2720 -648 2733 -644
rect 2737 -648 2740 -644
rect 3545 -645 3550 -643
rect 2713 -650 2740 -648
rect 3510 -650 3550 -645
rect 2721 -655 2725 -650
rect 3510 -654 3516 -653
rect 2219 -661 2246 -658
rect 2219 -665 2222 -661
rect 2226 -665 2239 -661
rect 2243 -665 2246 -661
rect 2219 -667 2246 -665
rect 2227 -672 2231 -667
rect 3510 -658 3511 -654
rect 3515 -658 3516 -654
rect 3510 -661 3516 -658
rect 3545 -661 3550 -650
rect 3605 -656 3614 -653
rect 3605 -660 3607 -656
rect 3611 -660 3614 -656
rect 3628 -660 3641 -657
rect 3605 -661 3614 -660
rect 3510 -665 3522 -661
rect 3510 -675 3516 -665
rect 3600 -665 3614 -661
rect 3542 -673 3560 -669
rect 3605 -673 3614 -665
rect 3510 -679 3511 -675
rect 3515 -679 3516 -675
rect 3510 -680 3516 -679
rect 3545 -683 3550 -673
rect 3605 -677 3607 -673
rect 3611 -677 3614 -673
rect 3605 -680 3614 -677
rect 3620 -683 3624 -680
rect 3574 -687 3624 -683
rect 3574 -692 3578 -687
rect 3510 -697 3578 -692
rect 3628 -693 3632 -680
rect 3635 -687 3641 -660
rect 3664 -687 3668 -677
rect 3635 -692 3656 -687
rect 3664 -692 3675 -687
rect 3510 -705 3516 -704
rect 3510 -709 3511 -705
rect 3515 -709 3516 -705
rect 3510 -712 3516 -709
rect 3545 -712 3550 -697
rect 3605 -707 3614 -704
rect 3605 -711 3607 -707
rect 3611 -711 3614 -707
rect 3605 -712 3614 -711
rect 3510 -716 3522 -712
rect 3510 -726 3516 -716
rect 3600 -716 3614 -712
rect 3542 -724 3560 -720
rect 3605 -724 3614 -716
rect 3510 -730 3511 -726
rect 3515 -730 3516 -726
rect 3510 -731 3516 -730
rect 2704 -743 2721 -738
rect 2729 -747 2733 -735
rect 3545 -744 3550 -724
rect 3605 -728 3607 -724
rect 3611 -728 3614 -724
rect 3605 -731 3614 -728
rect 3664 -695 3668 -692
rect 3620 -744 3624 -713
rect 3656 -721 3660 -715
rect 3648 -722 3675 -721
rect 3648 -726 3649 -722
rect 3653 -726 3670 -722
rect 3674 -726 3675 -722
rect 3648 -727 3675 -726
rect 3545 -747 3624 -744
rect 2210 -760 2227 -755
rect 2235 -764 2239 -752
rect 2227 -768 2239 -764
rect 2721 -751 2733 -747
rect 2721 -755 2725 -751
rect 2227 -772 2231 -768
rect 161 -797 188 -794
rect 161 -801 164 -797
rect 168 -801 181 -797
rect 185 -801 188 -797
rect 161 -803 188 -801
rect 169 -808 173 -803
rect 58 -816 63 -814
rect -74 -821 63 -816
rect -37 -1111 -28 -821
rect 23 -825 29 -824
rect 23 -829 24 -825
rect 28 -829 29 -825
rect 23 -832 29 -829
rect 58 -832 63 -821
rect 118 -827 127 -824
rect 118 -831 120 -827
rect 124 -831 127 -827
rect 141 -831 154 -828
rect 118 -832 127 -831
rect 23 -836 35 -832
rect 23 -846 29 -836
rect 113 -836 127 -832
rect 55 -844 73 -840
rect 118 -844 127 -836
rect 23 -850 24 -846
rect 28 -850 29 -846
rect 23 -851 29 -850
rect 58 -854 63 -844
rect 118 -848 120 -844
rect 124 -848 127 -844
rect 118 -851 127 -848
rect 133 -854 137 -851
rect 87 -858 137 -854
rect 87 -863 91 -858
rect -3 -868 91 -863
rect 141 -864 145 -851
rect 148 -858 154 -831
rect 177 -858 181 -848
rect 659 -850 713 -847
rect 659 -854 662 -850
rect 666 -854 679 -850
rect 683 -854 689 -850
rect 693 -854 706 -850
rect 710 -854 713 -850
rect 1377 -848 1431 -845
rect 1377 -852 1380 -848
rect 1384 -852 1397 -848
rect 1401 -852 1407 -848
rect 1411 -852 1424 -848
rect 1428 -852 1431 -848
rect 2268 -798 2295 -795
rect 2268 -802 2271 -798
rect 2275 -802 2288 -798
rect 2292 -802 2295 -798
rect 2268 -804 2295 -802
rect 2276 -809 2280 -804
rect 2762 -781 2789 -778
rect 2762 -785 2765 -781
rect 2769 -785 2782 -781
rect 2786 -785 2789 -781
rect 2762 -787 2789 -785
rect 2770 -792 2774 -787
rect 2697 -846 2706 -841
rect 2729 -842 2733 -835
rect 2778 -842 2782 -832
rect 1377 -854 1431 -852
rect 659 -856 713 -854
rect 148 -863 169 -858
rect 177 -863 188 -858
rect 667 -861 671 -856
rect 694 -861 698 -856
rect 997 -859 1051 -856
rect -12 -1045 -3 -868
rect 23 -876 29 -875
rect 23 -880 24 -876
rect 28 -880 29 -876
rect 23 -883 29 -880
rect 58 -883 63 -868
rect 118 -878 127 -875
rect 118 -882 120 -878
rect 124 -882 127 -878
rect 118 -883 127 -882
rect 23 -887 35 -883
rect 23 -897 29 -887
rect 113 -887 127 -883
rect 55 -895 73 -891
rect 118 -895 127 -887
rect 23 -901 24 -897
rect 28 -901 29 -897
rect 23 -902 29 -901
rect 58 -915 63 -895
rect 118 -899 120 -895
rect 124 -899 127 -895
rect 118 -902 127 -899
rect 177 -866 181 -863
rect 133 -915 137 -884
rect 169 -892 173 -886
rect 161 -893 188 -892
rect 161 -897 162 -893
rect 166 -897 183 -893
rect 187 -897 188 -893
rect 161 -898 188 -897
rect 997 -863 1000 -859
rect 1004 -863 1017 -859
rect 1021 -863 1027 -859
rect 1031 -863 1044 -859
rect 1048 -863 1051 -859
rect 997 -865 1051 -863
rect 1385 -859 1389 -854
rect 1412 -859 1416 -854
rect 58 -918 137 -915
rect 675 -921 679 -901
rect 702 -921 706 -901
rect 1005 -870 1009 -865
rect 1032 -870 1036 -865
rect 2203 -863 2212 -858
rect 2235 -859 2239 -852
rect 2284 -859 2288 -849
rect 2729 -847 2770 -842
rect 2778 -847 2789 -842
rect 2729 -850 2733 -847
rect 2778 -850 2782 -847
rect 2714 -854 2751 -850
rect 2235 -864 2276 -859
rect 2284 -864 2295 -859
rect 2714 -860 2718 -854
rect 2747 -860 2751 -854
rect 2235 -867 2239 -864
rect 2284 -867 2288 -864
rect 2220 -871 2257 -867
rect 2220 -877 2224 -871
rect 2253 -877 2257 -871
rect 721 -920 748 -917
rect 675 -925 716 -921
rect 660 -931 667 -926
rect 694 -935 698 -925
rect 58 -969 112 -966
rect 58 -973 61 -969
rect 65 -973 78 -969
rect 82 -973 88 -969
rect 92 -973 105 -969
rect 109 -973 112 -969
rect 58 -975 112 -973
rect 66 -980 70 -975
rect 93 -980 97 -975
rect 686 -981 690 -975
rect 711 -981 716 -925
rect 721 -924 724 -920
rect 728 -924 741 -920
rect 745 -924 748 -920
rect 721 -926 748 -924
rect 729 -931 733 -926
rect 1013 -930 1017 -910
rect 1040 -930 1044 -910
rect 1393 -919 1397 -899
rect 1420 -919 1424 -899
rect 2770 -876 2774 -870
rect 2762 -877 2789 -876
rect 2706 -886 2710 -880
rect 2739 -886 2743 -880
rect 2762 -881 2763 -877
rect 2767 -881 2784 -877
rect 2788 -881 2789 -877
rect 2762 -882 2789 -881
rect 2698 -887 2725 -886
rect 2276 -893 2280 -887
rect 2698 -891 2699 -887
rect 2703 -891 2720 -887
rect 2724 -891 2725 -887
rect 2698 -892 2725 -891
rect 2731 -887 2758 -886
rect 2731 -891 2732 -887
rect 2736 -891 2753 -887
rect 2757 -891 2758 -887
rect 2731 -892 2758 -891
rect 2268 -894 2295 -893
rect 2212 -903 2216 -897
rect 2245 -903 2249 -897
rect 2268 -898 2269 -894
rect 2273 -898 2290 -894
rect 2294 -898 2295 -894
rect 2268 -899 2295 -898
rect 2204 -904 2231 -903
rect 2204 -908 2205 -904
rect 2209 -908 2226 -904
rect 2230 -908 2231 -904
rect 2204 -909 2231 -908
rect 2237 -904 2264 -903
rect 2237 -908 2238 -904
rect 2242 -908 2259 -904
rect 2263 -908 2264 -904
rect 2237 -909 2264 -908
rect 1439 -918 1466 -915
rect 1393 -923 1434 -919
rect 1059 -929 1086 -926
rect 1378 -929 1385 -924
rect 1013 -934 1054 -930
rect 998 -940 1005 -935
rect 1032 -944 1036 -934
rect 737 -981 741 -971
rect 686 -985 700 -981
rect 694 -986 700 -985
rect 711 -986 729 -981
rect 737 -986 750 -981
rect 660 -997 686 -992
rect 694 -1000 698 -986
rect 737 -989 741 -986
rect 74 -1040 78 -1020
rect 101 -1040 105 -1020
rect 120 -1039 147 -1036
rect 74 -1044 115 -1040
rect -12 -1050 66 -1045
rect -12 -1051 -3 -1050
rect 93 -1054 97 -1044
rect 85 -1100 89 -1094
rect 110 -1100 115 -1044
rect 120 -1043 123 -1039
rect 127 -1043 140 -1039
rect 144 -1043 147 -1039
rect 120 -1045 147 -1043
rect 1024 -990 1028 -984
rect 1049 -990 1054 -934
rect 1059 -933 1062 -929
rect 1066 -933 1079 -929
rect 1083 -933 1086 -929
rect 1412 -933 1416 -923
rect 1059 -935 1086 -933
rect 1067 -940 1071 -935
rect 1075 -990 1079 -980
rect 1404 -979 1408 -973
rect 1429 -979 1434 -923
rect 1439 -922 1442 -918
rect 1446 -922 1459 -918
rect 1463 -922 1466 -918
rect 1439 -924 1466 -922
rect 1447 -929 1451 -924
rect 1455 -979 1459 -969
rect 1404 -983 1418 -979
rect 1412 -984 1418 -983
rect 1429 -984 1447 -979
rect 1455 -984 1468 -979
rect 1024 -994 1038 -990
rect 1032 -995 1038 -994
rect 1049 -995 1067 -990
rect 1075 -995 1088 -990
rect 1378 -995 1404 -990
rect 998 -1006 1024 -1001
rect 1032 -1009 1036 -995
rect 1075 -998 1079 -995
rect 1412 -998 1416 -984
rect 1455 -987 1459 -984
rect 729 -1015 733 -1009
rect 721 -1016 748 -1015
rect 721 -1020 722 -1016
rect 726 -1020 743 -1016
rect 747 -1020 748 -1016
rect 721 -1021 748 -1020
rect 128 -1050 132 -1045
rect 686 -1046 690 -1040
rect 678 -1047 705 -1046
rect 678 -1051 679 -1047
rect 683 -1051 700 -1047
rect 704 -1051 705 -1047
rect 678 -1052 705 -1051
rect 1067 -1024 1071 -1018
rect 1059 -1025 1086 -1024
rect 1059 -1029 1060 -1025
rect 1064 -1029 1081 -1025
rect 1085 -1029 1086 -1025
rect 1059 -1030 1086 -1029
rect 1447 -1013 1451 -1007
rect 1439 -1014 1466 -1013
rect 1439 -1018 1440 -1014
rect 1444 -1018 1461 -1014
rect 1465 -1018 1466 -1014
rect 1439 -1019 1466 -1018
rect 1404 -1044 1408 -1038
rect 1396 -1045 1423 -1044
rect 1396 -1049 1397 -1045
rect 1401 -1049 1418 -1045
rect 1422 -1049 1423 -1045
rect 1024 -1055 1028 -1049
rect 1396 -1050 1423 -1049
rect 1016 -1056 1043 -1055
rect 1016 -1060 1017 -1056
rect 1021 -1060 1038 -1056
rect 1042 -1060 1043 -1056
rect 1016 -1061 1043 -1060
rect 136 -1100 140 -1090
rect 85 -1104 99 -1100
rect 93 -1105 99 -1104
rect 110 -1105 128 -1100
rect 136 -1105 149 -1100
rect -37 -1116 85 -1111
rect 93 -1119 97 -1105
rect 136 -1108 140 -1105
rect 128 -1134 132 -1128
rect 120 -1135 147 -1134
rect 120 -1139 121 -1135
rect 125 -1139 142 -1135
rect 146 -1139 147 -1135
rect 120 -1140 147 -1139
rect 85 -1165 89 -1159
rect 77 -1166 104 -1165
rect 77 -1170 78 -1166
rect 82 -1170 99 -1166
rect 103 -1170 104 -1166
rect 77 -1171 104 -1170
rect 5974 -1721 6001 -1718
rect 5974 -1725 5977 -1721
rect 5981 -1725 5994 -1721
rect 5998 -1725 6001 -1721
rect 5974 -1727 6001 -1725
rect 5982 -1732 5986 -1727
rect 5871 -1740 5876 -1738
rect 5836 -1745 5876 -1740
rect 5836 -1749 5842 -1748
rect 5836 -1753 5837 -1749
rect 5841 -1753 5842 -1749
rect 5836 -1756 5842 -1753
rect 5871 -1756 5876 -1745
rect 5931 -1751 5940 -1748
rect 5931 -1755 5933 -1751
rect 5937 -1755 5940 -1751
rect 5954 -1755 5967 -1752
rect 5931 -1756 5940 -1755
rect 4921 -1762 4948 -1759
rect 4002 -1768 4029 -1765
rect 4921 -1766 4924 -1762
rect 4928 -1766 4941 -1762
rect 4945 -1766 4948 -1762
rect 4921 -1768 4948 -1766
rect 5836 -1760 5848 -1756
rect 4002 -1772 4005 -1768
rect 4009 -1772 4022 -1768
rect 4026 -1772 4029 -1768
rect 4002 -1774 4029 -1772
rect 4929 -1773 4933 -1768
rect 5836 -1770 5842 -1760
rect 5926 -1760 5940 -1756
rect 5868 -1768 5886 -1764
rect 5931 -1768 5940 -1760
rect 4010 -1779 4014 -1774
rect 4456 -1797 4483 -1794
rect 4456 -1801 4459 -1797
rect 4463 -1801 4476 -1797
rect 4480 -1801 4483 -1797
rect 4456 -1803 4483 -1801
rect 2164 -1864 2218 -1861
rect 2164 -1868 2167 -1864
rect 2171 -1868 2184 -1864
rect 2188 -1868 2194 -1864
rect 2198 -1868 2211 -1864
rect 2215 -1868 2218 -1864
rect 2164 -1870 2218 -1868
rect 2769 -1864 2823 -1861
rect 2769 -1868 2772 -1864
rect 2776 -1868 2789 -1864
rect 2793 -1868 2799 -1864
rect 2803 -1868 2816 -1864
rect 2820 -1868 2823 -1864
rect 2769 -1870 2823 -1868
rect 3374 -1864 3428 -1861
rect 3374 -1868 3377 -1864
rect 3381 -1868 3394 -1864
rect 3398 -1868 3404 -1864
rect 3408 -1868 3421 -1864
rect 3425 -1868 3428 -1864
rect 3993 -1867 4010 -1862
rect 3374 -1870 3428 -1868
rect 2172 -1875 2176 -1870
rect 2199 -1875 2203 -1870
rect 2777 -1875 2781 -1870
rect 2804 -1875 2808 -1870
rect 3382 -1875 3386 -1870
rect 3409 -1875 3413 -1870
rect 4018 -1871 4022 -1859
rect 4010 -1875 4022 -1871
rect 4464 -1808 4468 -1803
rect 1663 -1899 1717 -1896
rect 1261 -1902 1315 -1899
rect 1261 -1906 1264 -1902
rect 1268 -1906 1281 -1902
rect 1285 -1906 1291 -1902
rect 1295 -1906 1308 -1902
rect 1312 -1906 1315 -1902
rect 1663 -1903 1666 -1899
rect 1670 -1903 1683 -1899
rect 1687 -1903 1693 -1899
rect 1697 -1903 1710 -1899
rect 1714 -1903 1717 -1899
rect 1663 -1905 1717 -1903
rect 1261 -1908 1315 -1906
rect 793 -1911 847 -1908
rect 793 -1915 796 -1911
rect 800 -1915 813 -1911
rect 817 -1915 823 -1911
rect 827 -1915 840 -1911
rect 844 -1915 847 -1911
rect 793 -1917 847 -1915
rect 1269 -1913 1273 -1908
rect 1296 -1913 1300 -1908
rect 1671 -1910 1675 -1905
rect 1698 -1910 1702 -1905
rect 146 -1921 173 -1918
rect 146 -1925 149 -1921
rect 153 -1925 166 -1921
rect 170 -1925 173 -1921
rect 146 -1927 173 -1925
rect 801 -1922 805 -1917
rect 828 -1922 832 -1917
rect 154 -1932 158 -1927
rect 43 -1940 48 -1938
rect -89 -1945 48 -1940
rect -52 -2235 -43 -1945
rect 8 -1949 14 -1948
rect 8 -1953 9 -1949
rect 13 -1953 14 -1949
rect 8 -1956 14 -1953
rect 43 -1956 48 -1945
rect 103 -1951 112 -1948
rect 103 -1955 105 -1951
rect 109 -1955 112 -1951
rect 126 -1955 139 -1952
rect 103 -1956 112 -1955
rect 8 -1960 20 -1956
rect 8 -1970 14 -1960
rect 98 -1960 112 -1956
rect 40 -1968 58 -1964
rect 103 -1968 112 -1960
rect 8 -1974 9 -1970
rect 13 -1974 14 -1970
rect 8 -1975 14 -1974
rect 43 -1978 48 -1968
rect 103 -1972 105 -1968
rect 109 -1972 112 -1968
rect 103 -1975 112 -1972
rect 118 -1978 122 -1975
rect 72 -1982 122 -1978
rect 72 -1987 76 -1982
rect -18 -1992 76 -1987
rect 126 -1988 130 -1975
rect 133 -1982 139 -1955
rect 2180 -1935 2184 -1915
rect 2207 -1935 2211 -1915
rect 2226 -1934 2253 -1931
rect 2180 -1939 2221 -1935
rect 2165 -1945 2172 -1940
rect 2199 -1949 2203 -1939
rect 162 -1982 166 -1972
rect 809 -1982 813 -1962
rect 836 -1982 840 -1962
rect 1277 -1973 1281 -1953
rect 1304 -1973 1308 -1953
rect 1323 -1972 1350 -1969
rect 1277 -1977 1318 -1973
rect 855 -1981 882 -1978
rect 133 -1987 154 -1982
rect 162 -1987 173 -1982
rect 809 -1986 850 -1982
rect -27 -2169 -18 -1992
rect 8 -2000 14 -1999
rect 8 -2004 9 -2000
rect 13 -2004 14 -2000
rect 8 -2007 14 -2004
rect 43 -2007 48 -1992
rect 103 -2002 112 -1999
rect 103 -2006 105 -2002
rect 109 -2006 112 -2002
rect 103 -2007 112 -2006
rect 8 -2011 20 -2007
rect 8 -2021 14 -2011
rect 98 -2011 112 -2007
rect 40 -2019 58 -2015
rect 103 -2019 112 -2011
rect 8 -2025 9 -2021
rect 13 -2025 14 -2021
rect 8 -2026 14 -2025
rect 43 -2039 48 -2019
rect 103 -2023 105 -2019
rect 109 -2023 112 -2019
rect 103 -2026 112 -2023
rect 162 -1990 166 -1987
rect 118 -2039 122 -2008
rect 794 -1992 801 -1987
rect 828 -1996 832 -1986
rect 154 -2016 158 -2010
rect 146 -2017 173 -2016
rect 146 -2021 147 -2017
rect 151 -2021 168 -2017
rect 172 -2021 173 -2017
rect 146 -2022 173 -2021
rect 43 -2042 122 -2039
rect 820 -2042 824 -2036
rect 845 -2042 850 -1986
rect 855 -1985 858 -1981
rect 862 -1985 875 -1981
rect 879 -1985 882 -1981
rect 1262 -1983 1269 -1978
rect 855 -1987 882 -1985
rect 1296 -1987 1300 -1977
rect 863 -1992 867 -1987
rect 871 -2042 875 -2032
rect 1288 -2033 1292 -2027
rect 1313 -2033 1318 -1977
rect 1323 -1976 1326 -1972
rect 1330 -1976 1343 -1972
rect 1347 -1976 1350 -1972
rect 1679 -1970 1683 -1950
rect 1706 -1970 1710 -1950
rect 1725 -1969 1752 -1966
rect 1679 -1974 1720 -1970
rect 1323 -1978 1350 -1976
rect 1331 -1983 1335 -1978
rect 1664 -1980 1671 -1975
rect 1698 -1984 1702 -1974
rect 1339 -2033 1343 -2023
rect 1690 -2030 1694 -2024
rect 1715 -2030 1720 -1974
rect 1725 -1973 1728 -1969
rect 1732 -1973 1745 -1969
rect 1749 -1973 1752 -1969
rect 1725 -1975 1752 -1973
rect 1733 -1980 1737 -1975
rect 2191 -1995 2195 -1989
rect 2216 -1995 2221 -1939
rect 2226 -1938 2229 -1934
rect 2233 -1938 2246 -1934
rect 2250 -1938 2253 -1934
rect 2226 -1940 2253 -1938
rect 2785 -1935 2789 -1915
rect 2812 -1935 2816 -1915
rect 2831 -1934 2858 -1931
rect 2785 -1939 2826 -1935
rect 2234 -1945 2238 -1940
rect 2770 -1945 2777 -1940
rect 2804 -1949 2808 -1939
rect 2242 -1995 2246 -1985
rect 2796 -1995 2800 -1989
rect 2821 -1995 2826 -1939
rect 2831 -1938 2834 -1934
rect 2838 -1938 2851 -1934
rect 2855 -1938 2858 -1934
rect 2831 -1940 2858 -1938
rect 3390 -1935 3394 -1915
rect 3417 -1935 3421 -1915
rect 4010 -1879 4014 -1875
rect 3436 -1934 3463 -1931
rect 3390 -1939 3431 -1935
rect 2839 -1945 2843 -1940
rect 3375 -1945 3382 -1940
rect 3409 -1949 3413 -1939
rect 2847 -1995 2851 -1985
rect 3401 -1995 3405 -1989
rect 3426 -1995 3431 -1939
rect 3436 -1938 3439 -1934
rect 3443 -1938 3456 -1934
rect 3460 -1938 3463 -1934
rect 3436 -1940 3463 -1938
rect 3444 -1945 3448 -1940
rect 5836 -1774 5837 -1770
rect 5841 -1774 5842 -1770
rect 5836 -1775 5842 -1774
rect 5871 -1778 5876 -1768
rect 5931 -1772 5933 -1768
rect 5937 -1772 5940 -1768
rect 5931 -1775 5940 -1772
rect 5946 -1778 5950 -1775
rect 5900 -1782 5950 -1778
rect 5900 -1787 5904 -1782
rect 5836 -1792 5904 -1787
rect 5954 -1788 5958 -1775
rect 5961 -1782 5967 -1755
rect 5990 -1782 5994 -1772
rect 5961 -1787 5982 -1782
rect 5990 -1787 6001 -1782
rect 5836 -1800 5842 -1799
rect 5836 -1804 5837 -1800
rect 5841 -1804 5842 -1800
rect 5836 -1807 5842 -1804
rect 5871 -1807 5876 -1792
rect 5931 -1802 5940 -1799
rect 5931 -1806 5933 -1802
rect 5937 -1806 5940 -1802
rect 5931 -1807 5940 -1806
rect 5836 -1811 5848 -1807
rect 5836 -1821 5842 -1811
rect 5926 -1811 5940 -1807
rect 5868 -1819 5886 -1815
rect 5931 -1819 5940 -1811
rect 5836 -1825 5837 -1821
rect 5841 -1825 5842 -1821
rect 5836 -1826 5842 -1825
rect 5871 -1839 5876 -1819
rect 5931 -1823 5933 -1819
rect 5937 -1823 5940 -1819
rect 5931 -1826 5940 -1823
rect 5990 -1790 5994 -1787
rect 5946 -1839 5950 -1808
rect 5982 -1816 5986 -1810
rect 5974 -1817 6001 -1816
rect 5974 -1821 5975 -1817
rect 5979 -1821 5996 -1817
rect 6000 -1821 6001 -1817
rect 5974 -1822 6001 -1821
rect 5871 -1842 5950 -1839
rect 4912 -1861 4929 -1856
rect 4937 -1865 4941 -1853
rect 4447 -1896 4464 -1891
rect 4472 -1900 4476 -1888
rect 4051 -1905 4078 -1902
rect 4051 -1909 4054 -1905
rect 4058 -1909 4071 -1905
rect 4075 -1909 4078 -1905
rect 4051 -1911 4078 -1909
rect 4464 -1904 4476 -1900
rect 4929 -1869 4941 -1865
rect 4929 -1873 4933 -1869
rect 4464 -1908 4468 -1904
rect 4059 -1916 4063 -1911
rect 3986 -1970 3995 -1965
rect 4018 -1966 4022 -1959
rect 4067 -1966 4071 -1956
rect 4018 -1971 4059 -1966
rect 4067 -1971 4078 -1966
rect 4018 -1974 4022 -1971
rect 4067 -1974 4071 -1971
rect 4003 -1978 4040 -1974
rect 4003 -1984 4007 -1978
rect 4036 -1984 4040 -1978
rect 3452 -1995 3456 -1985
rect 2191 -1999 2205 -1995
rect 2199 -2000 2205 -1999
rect 2216 -2000 2234 -1995
rect 2242 -2000 2255 -1995
rect 2796 -1999 2810 -1995
rect 2804 -2000 2810 -1999
rect 2821 -2000 2839 -1995
rect 2847 -2000 2860 -1995
rect 3401 -1999 3415 -1995
rect 3409 -2000 3415 -1999
rect 3426 -2000 3444 -1995
rect 3452 -2000 3465 -1995
rect 2165 -2011 2191 -2006
rect 2199 -2014 2203 -2000
rect 2242 -2003 2246 -2000
rect 1741 -2030 1745 -2020
rect 1288 -2037 1302 -2033
rect 1296 -2038 1302 -2037
rect 1313 -2038 1331 -2033
rect 1339 -2038 1352 -2033
rect 1690 -2034 1704 -2030
rect 1698 -2035 1704 -2034
rect 1715 -2035 1733 -2030
rect 1741 -2035 1754 -2030
rect 820 -2046 834 -2042
rect 828 -2047 834 -2046
rect 845 -2047 863 -2042
rect 871 -2047 884 -2042
rect 794 -2058 820 -2053
rect 828 -2061 832 -2047
rect 871 -2050 875 -2047
rect 1262 -2049 1288 -2044
rect 43 -2093 97 -2090
rect 43 -2097 46 -2093
rect 50 -2097 63 -2093
rect 67 -2097 73 -2093
rect 77 -2097 90 -2093
rect 94 -2097 97 -2093
rect 43 -2099 97 -2097
rect 51 -2104 55 -2099
rect 78 -2104 82 -2099
rect 1296 -2052 1300 -2038
rect 1339 -2041 1343 -2038
rect 863 -2076 867 -2070
rect 855 -2077 882 -2076
rect 855 -2081 856 -2077
rect 860 -2081 877 -2077
rect 881 -2081 882 -2077
rect 855 -2082 882 -2081
rect 1664 -2046 1690 -2041
rect 1698 -2049 1702 -2035
rect 1741 -2038 1745 -2035
rect 1331 -2067 1335 -2061
rect 1323 -2068 1350 -2067
rect 1323 -2072 1324 -2068
rect 1328 -2072 1345 -2068
rect 1349 -2072 1350 -2068
rect 1323 -2073 1350 -2072
rect 2770 -2011 2796 -2006
rect 2804 -2014 2808 -2000
rect 2847 -2003 2851 -2000
rect 2234 -2029 2238 -2023
rect 2226 -2030 2253 -2029
rect 2226 -2034 2227 -2030
rect 2231 -2034 2248 -2030
rect 2252 -2034 2253 -2030
rect 2226 -2035 2253 -2034
rect 3375 -2011 3401 -2006
rect 3409 -2014 3413 -2000
rect 3452 -2003 3456 -2000
rect 2839 -2029 2843 -2023
rect 2831 -2030 2858 -2029
rect 2831 -2034 2832 -2030
rect 2836 -2034 2853 -2030
rect 2857 -2034 2858 -2030
rect 2831 -2035 2858 -2034
rect 4505 -1934 4532 -1931
rect 4505 -1938 4508 -1934
rect 4512 -1938 4525 -1934
rect 4529 -1938 4532 -1934
rect 4505 -1940 4532 -1938
rect 4513 -1945 4517 -1940
rect 4970 -1899 4997 -1896
rect 4970 -1903 4973 -1899
rect 4977 -1903 4990 -1899
rect 4994 -1903 4997 -1899
rect 4970 -1905 4997 -1903
rect 4978 -1910 4982 -1905
rect 4905 -1964 4914 -1959
rect 4937 -1960 4941 -1953
rect 4986 -1960 4990 -1950
rect 4937 -1965 4978 -1960
rect 4986 -1965 4997 -1960
rect 4937 -1968 4941 -1965
rect 4986 -1968 4990 -1965
rect 4922 -1972 4959 -1968
rect 4922 -1978 4926 -1972
rect 4955 -1978 4959 -1972
rect 4059 -2000 4063 -1994
rect 4440 -1999 4449 -1994
rect 4472 -1995 4476 -1988
rect 4521 -1995 4525 -1985
rect 4472 -2000 4513 -1995
rect 4521 -2000 4532 -1995
rect 4978 -1994 4982 -1988
rect 4970 -1995 4997 -1994
rect 4051 -2001 4078 -2000
rect 3995 -2010 3999 -2004
rect 4028 -2010 4032 -2004
rect 4051 -2005 4052 -2001
rect 4056 -2005 4073 -2001
rect 4077 -2005 4078 -2001
rect 4472 -2003 4476 -2000
rect 4521 -2003 4525 -2000
rect 4051 -2006 4078 -2005
rect 4457 -2007 4494 -2003
rect 3987 -2011 4014 -2010
rect 3987 -2015 3988 -2011
rect 3992 -2015 4009 -2011
rect 4013 -2015 4014 -2011
rect 3987 -2016 4014 -2015
rect 4020 -2011 4047 -2010
rect 4020 -2015 4021 -2011
rect 4025 -2015 4042 -2011
rect 4046 -2015 4047 -2011
rect 4457 -2013 4461 -2007
rect 4490 -2013 4494 -2007
rect 4020 -2016 4047 -2015
rect 3444 -2029 3448 -2023
rect 3436 -2030 3463 -2029
rect 3436 -2034 3437 -2030
rect 3441 -2034 3458 -2030
rect 3462 -2034 3463 -2030
rect 3436 -2035 3463 -2034
rect 4914 -2004 4918 -1998
rect 4947 -2004 4951 -1998
rect 4970 -1999 4971 -1995
rect 4975 -1999 4992 -1995
rect 4996 -1999 4997 -1995
rect 4970 -2000 4997 -1999
rect 4906 -2005 4933 -2004
rect 4906 -2009 4907 -2005
rect 4911 -2009 4928 -2005
rect 4932 -2009 4933 -2005
rect 4906 -2010 4933 -2009
rect 4939 -2005 4966 -2004
rect 4939 -2009 4940 -2005
rect 4944 -2009 4961 -2005
rect 4965 -2009 4966 -2005
rect 4939 -2010 4966 -2009
rect 4513 -2029 4517 -2023
rect 4505 -2030 4532 -2029
rect 4449 -2039 4453 -2033
rect 4482 -2039 4486 -2033
rect 4505 -2034 4506 -2030
rect 4510 -2034 4527 -2030
rect 4531 -2034 4532 -2030
rect 4505 -2035 4532 -2034
rect 4441 -2040 4468 -2039
rect 4441 -2044 4442 -2040
rect 4446 -2044 4463 -2040
rect 4467 -2044 4468 -2040
rect 4441 -2045 4468 -2044
rect 4474 -2040 4501 -2039
rect 4474 -2044 4475 -2040
rect 4479 -2044 4496 -2040
rect 4500 -2044 4501 -2040
rect 4474 -2045 4501 -2044
rect 1733 -2064 1737 -2058
rect 2191 -2060 2195 -2054
rect 2796 -2060 2800 -2054
rect 3401 -2060 3405 -2054
rect 2183 -2061 2210 -2060
rect 1725 -2065 1752 -2064
rect 1725 -2069 1726 -2065
rect 1730 -2069 1747 -2065
rect 1751 -2069 1752 -2065
rect 2183 -2065 2184 -2061
rect 2188 -2065 2205 -2061
rect 2209 -2065 2210 -2061
rect 2183 -2066 2210 -2065
rect 2788 -2061 2815 -2060
rect 2788 -2065 2789 -2061
rect 2793 -2065 2810 -2061
rect 2814 -2065 2815 -2061
rect 2788 -2066 2815 -2065
rect 3393 -2061 3420 -2060
rect 3393 -2065 3394 -2061
rect 3398 -2065 3415 -2061
rect 3419 -2065 3420 -2061
rect 3393 -2066 3420 -2065
rect 1725 -2070 1752 -2069
rect 1288 -2098 1292 -2092
rect 1690 -2095 1694 -2089
rect 1682 -2096 1709 -2095
rect 1280 -2099 1307 -2098
rect 820 -2107 824 -2101
rect 1280 -2103 1281 -2099
rect 1285 -2103 1302 -2099
rect 1306 -2103 1307 -2099
rect 1682 -2100 1683 -2096
rect 1687 -2100 1704 -2096
rect 1708 -2100 1709 -2096
rect 1682 -2101 1709 -2100
rect 1280 -2104 1307 -2103
rect 812 -2108 839 -2107
rect 812 -2112 813 -2108
rect 817 -2112 834 -2108
rect 838 -2112 839 -2108
rect 812 -2113 839 -2112
rect 59 -2164 63 -2144
rect 86 -2164 90 -2144
rect 105 -2163 132 -2160
rect 59 -2168 100 -2164
rect -27 -2174 51 -2169
rect -27 -2175 -18 -2174
rect 78 -2178 82 -2168
rect 70 -2224 74 -2218
rect 95 -2224 100 -2168
rect 105 -2167 108 -2163
rect 112 -2167 125 -2163
rect 129 -2167 132 -2163
rect 105 -2169 132 -2167
rect 113 -2174 117 -2169
rect 121 -2224 125 -2214
rect 70 -2228 84 -2224
rect 78 -2229 84 -2228
rect 95 -2229 113 -2224
rect 121 -2229 134 -2224
rect -52 -2240 70 -2235
rect 78 -2243 82 -2229
rect 121 -2232 125 -2229
rect 113 -2258 117 -2252
rect 105 -2259 132 -2258
rect 105 -2263 106 -2259
rect 110 -2263 127 -2259
rect 131 -2263 132 -2259
rect 105 -2264 132 -2263
rect 70 -2289 74 -2283
rect 62 -2290 89 -2289
rect 62 -2294 63 -2290
rect 67 -2294 84 -2290
rect 88 -2294 89 -2290
rect 62 -2295 89 -2294
rect 7407 -3113 7434 -3110
rect 6488 -3119 6515 -3116
rect 7407 -3117 7410 -3113
rect 7414 -3117 7427 -3113
rect 7431 -3117 7434 -3113
rect 7407 -3119 7434 -3117
rect 6057 -3125 6084 -3122
rect 6488 -3123 6491 -3119
rect 6495 -3123 6508 -3119
rect 6512 -3123 6515 -3119
rect 6488 -3125 6515 -3123
rect 7415 -3124 7419 -3119
rect 6057 -3129 6060 -3125
rect 6064 -3129 6077 -3125
rect 6081 -3129 6084 -3125
rect 6057 -3131 6084 -3129
rect 6496 -3130 6500 -3125
rect 6065 -3136 6069 -3131
rect 6942 -3148 6969 -3145
rect 6942 -3152 6945 -3148
rect 6949 -3152 6962 -3148
rect 6966 -3152 6969 -3148
rect 6942 -3154 6969 -3152
rect 6048 -3224 6065 -3219
rect 6073 -3228 6077 -3216
rect 6479 -3218 6496 -3213
rect 6504 -3222 6508 -3210
rect 6065 -3232 6077 -3228
rect 6496 -3226 6508 -3222
rect 6950 -3159 6954 -3154
rect 6496 -3230 6500 -3226
rect 6065 -3236 6069 -3232
rect 4204 -3289 4258 -3286
rect 4204 -3293 4207 -3289
rect 4211 -3293 4224 -3289
rect 4228 -3293 4234 -3289
rect 4238 -3293 4251 -3289
rect 4255 -3293 4258 -3289
rect 4204 -3295 4258 -3293
rect 4212 -3300 4216 -3295
rect 4239 -3300 4243 -3295
rect 2711 -3306 2765 -3303
rect 2711 -3310 2714 -3306
rect 2718 -3310 2731 -3306
rect 2735 -3310 2741 -3306
rect 2745 -3310 2758 -3306
rect 2762 -3310 2765 -3306
rect 3429 -3304 3483 -3301
rect 3429 -3308 3432 -3304
rect 3436 -3308 3449 -3304
rect 3453 -3308 3459 -3304
rect 3463 -3308 3476 -3304
rect 3480 -3308 3483 -3304
rect 3429 -3310 3483 -3308
rect 2711 -3312 2765 -3310
rect 2719 -3317 2723 -3312
rect 2746 -3317 2750 -3312
rect 3049 -3315 3103 -3312
rect 884 -3337 938 -3334
rect 146 -3340 173 -3337
rect 146 -3344 149 -3340
rect 153 -3344 166 -3340
rect 170 -3344 173 -3340
rect 884 -3341 887 -3337
rect 891 -3341 904 -3337
rect 908 -3341 914 -3337
rect 918 -3341 931 -3337
rect 935 -3341 938 -3337
rect 1602 -3335 1656 -3332
rect 1602 -3339 1605 -3335
rect 1609 -3339 1622 -3335
rect 1626 -3339 1632 -3335
rect 1636 -3339 1649 -3335
rect 1653 -3339 1656 -3335
rect 1602 -3341 1656 -3339
rect 884 -3343 938 -3341
rect 146 -3346 173 -3344
rect 154 -3351 158 -3346
rect 892 -3348 896 -3343
rect 919 -3348 923 -3343
rect 1222 -3346 1276 -3343
rect 43 -3359 48 -3357
rect -89 -3364 48 -3359
rect -52 -3654 -43 -3364
rect 8 -3368 14 -3367
rect 8 -3372 9 -3368
rect 13 -3372 14 -3368
rect 8 -3375 14 -3372
rect 43 -3375 48 -3364
rect 103 -3370 112 -3367
rect 103 -3374 105 -3370
rect 109 -3374 112 -3370
rect 126 -3374 139 -3371
rect 103 -3375 112 -3374
rect 8 -3379 20 -3375
rect 8 -3389 14 -3379
rect 98 -3379 112 -3375
rect 40 -3387 58 -3383
rect 103 -3387 112 -3379
rect 8 -3393 9 -3389
rect 13 -3393 14 -3389
rect 8 -3394 14 -3393
rect 43 -3397 48 -3387
rect 103 -3391 105 -3387
rect 109 -3391 112 -3387
rect 103 -3394 112 -3391
rect 118 -3397 122 -3394
rect 72 -3401 122 -3397
rect 72 -3406 76 -3401
rect -18 -3411 76 -3406
rect 126 -3407 130 -3394
rect 133 -3401 139 -3374
rect 1222 -3350 1225 -3346
rect 1229 -3350 1242 -3346
rect 1246 -3350 1252 -3346
rect 1256 -3350 1269 -3346
rect 1273 -3350 1276 -3346
rect 1222 -3352 1276 -3350
rect 1610 -3346 1614 -3341
rect 1637 -3346 1641 -3341
rect 162 -3401 166 -3391
rect 133 -3406 154 -3401
rect 162 -3406 173 -3401
rect -27 -3588 -18 -3411
rect 8 -3419 14 -3418
rect 8 -3423 9 -3419
rect 13 -3423 14 -3419
rect 8 -3426 14 -3423
rect 43 -3426 48 -3411
rect 103 -3421 112 -3418
rect 103 -3425 105 -3421
rect 109 -3425 112 -3421
rect 103 -3426 112 -3425
rect 8 -3430 20 -3426
rect 8 -3440 14 -3430
rect 98 -3430 112 -3426
rect 40 -3438 58 -3434
rect 103 -3438 112 -3430
rect 8 -3444 9 -3440
rect 13 -3444 14 -3440
rect 8 -3445 14 -3444
rect 43 -3458 48 -3438
rect 103 -3442 105 -3438
rect 109 -3442 112 -3438
rect 103 -3445 112 -3442
rect 162 -3409 166 -3406
rect 118 -3458 122 -3427
rect 900 -3408 904 -3388
rect 927 -3408 931 -3388
rect 1230 -3357 1234 -3352
rect 1257 -3357 1261 -3352
rect 3049 -3319 3052 -3315
rect 3056 -3319 3069 -3315
rect 3073 -3319 3079 -3315
rect 3083 -3319 3096 -3315
rect 3100 -3319 3103 -3315
rect 3049 -3321 3103 -3319
rect 3437 -3315 3441 -3310
rect 3464 -3315 3468 -3310
rect 2727 -3377 2731 -3357
rect 2754 -3377 2758 -3357
rect 3057 -3326 3061 -3321
rect 3084 -3326 3088 -3321
rect 4526 -3303 4580 -3300
rect 4526 -3307 4529 -3303
rect 4533 -3307 4546 -3303
rect 4550 -3307 4556 -3303
rect 4560 -3307 4573 -3303
rect 4577 -3307 4580 -3303
rect 5244 -3301 5298 -3298
rect 5244 -3305 5247 -3301
rect 5251 -3305 5264 -3301
rect 5268 -3305 5274 -3301
rect 5278 -3305 5291 -3301
rect 5295 -3305 5298 -3301
rect 5244 -3307 5298 -3305
rect 4526 -3309 4580 -3307
rect 2773 -3376 2800 -3373
rect 2727 -3381 2768 -3377
rect 946 -3407 973 -3404
rect 900 -3412 941 -3408
rect 885 -3418 892 -3413
rect 919 -3422 923 -3412
rect 154 -3435 158 -3429
rect 146 -3436 173 -3435
rect 146 -3440 147 -3436
rect 151 -3440 168 -3436
rect 172 -3440 173 -3436
rect 146 -3441 173 -3440
rect 43 -3461 122 -3458
rect 911 -3468 915 -3462
rect 936 -3468 941 -3412
rect 946 -3411 949 -3407
rect 953 -3411 966 -3407
rect 970 -3411 973 -3407
rect 946 -3413 973 -3411
rect 954 -3418 958 -3413
rect 1238 -3417 1242 -3397
rect 1265 -3417 1269 -3397
rect 1618 -3406 1622 -3386
rect 1645 -3406 1649 -3386
rect 2712 -3387 2719 -3382
rect 2746 -3391 2750 -3381
rect 1664 -3405 1691 -3402
rect 1618 -3410 1659 -3406
rect 1284 -3416 1311 -3413
rect 1603 -3416 1610 -3411
rect 1238 -3421 1279 -3417
rect 1223 -3427 1230 -3422
rect 1257 -3431 1261 -3421
rect 962 -3468 966 -3458
rect 911 -3472 925 -3468
rect 919 -3473 925 -3472
rect 936 -3473 954 -3468
rect 962 -3473 975 -3468
rect 885 -3484 911 -3479
rect 919 -3487 923 -3473
rect 962 -3476 966 -3473
rect 43 -3512 97 -3509
rect 43 -3516 46 -3512
rect 50 -3516 63 -3512
rect 67 -3516 73 -3512
rect 77 -3516 90 -3512
rect 94 -3516 97 -3512
rect 43 -3518 97 -3516
rect 51 -3523 55 -3518
rect 78 -3523 82 -3518
rect 1249 -3477 1253 -3471
rect 1274 -3477 1279 -3421
rect 1284 -3420 1287 -3416
rect 1291 -3420 1304 -3416
rect 1308 -3420 1311 -3416
rect 1637 -3420 1641 -3410
rect 1284 -3422 1311 -3420
rect 1292 -3427 1296 -3422
rect 1300 -3477 1304 -3467
rect 1629 -3466 1633 -3460
rect 1654 -3466 1659 -3410
rect 1664 -3409 1667 -3405
rect 1671 -3409 1684 -3405
rect 1688 -3409 1691 -3405
rect 1664 -3411 1691 -3409
rect 1672 -3416 1676 -3411
rect 2738 -3437 2742 -3431
rect 2763 -3437 2768 -3381
rect 2773 -3380 2776 -3376
rect 2780 -3380 2793 -3376
rect 2797 -3380 2800 -3376
rect 2773 -3382 2800 -3380
rect 2781 -3387 2785 -3382
rect 3065 -3386 3069 -3366
rect 3092 -3386 3096 -3366
rect 3445 -3375 3449 -3355
rect 3472 -3375 3476 -3355
rect 4220 -3360 4224 -3340
rect 4247 -3360 4251 -3340
rect 4534 -3314 4538 -3309
rect 4561 -3314 4565 -3309
rect 4864 -3312 4918 -3309
rect 4864 -3316 4867 -3312
rect 4871 -3316 4884 -3312
rect 4888 -3316 4894 -3312
rect 4898 -3316 4911 -3312
rect 4915 -3316 4918 -3312
rect 4864 -3318 4918 -3316
rect 5252 -3312 5256 -3307
rect 5279 -3312 5283 -3307
rect 4266 -3359 4293 -3356
rect 4220 -3364 4261 -3360
rect 4205 -3370 4212 -3365
rect 3491 -3374 3518 -3371
rect 4239 -3374 4243 -3364
rect 3445 -3379 3486 -3375
rect 3111 -3385 3138 -3382
rect 3430 -3385 3437 -3380
rect 3065 -3390 3106 -3386
rect 3050 -3396 3057 -3391
rect 3084 -3400 3088 -3390
rect 2789 -3437 2793 -3427
rect 2738 -3441 2752 -3437
rect 2746 -3442 2752 -3441
rect 2763 -3442 2781 -3437
rect 2789 -3442 2802 -3437
rect 2712 -3453 2738 -3448
rect 2746 -3456 2750 -3442
rect 2789 -3445 2793 -3442
rect 1680 -3466 1684 -3456
rect 1629 -3470 1643 -3466
rect 1637 -3471 1643 -3470
rect 1654 -3471 1672 -3466
rect 1680 -3471 1693 -3466
rect 1249 -3481 1263 -3477
rect 1257 -3482 1263 -3481
rect 1274 -3482 1292 -3477
rect 1300 -3482 1313 -3477
rect 1603 -3482 1629 -3477
rect 1223 -3493 1249 -3488
rect 1257 -3496 1261 -3482
rect 1300 -3485 1304 -3482
rect 1637 -3485 1641 -3471
rect 1680 -3474 1684 -3471
rect 954 -3502 958 -3496
rect 946 -3503 973 -3502
rect 946 -3507 947 -3503
rect 951 -3507 968 -3503
rect 972 -3507 973 -3503
rect 946 -3508 973 -3507
rect 911 -3533 915 -3527
rect 903 -3534 930 -3533
rect 903 -3538 904 -3534
rect 908 -3538 925 -3534
rect 929 -3538 930 -3534
rect 903 -3539 930 -3538
rect 1292 -3511 1296 -3505
rect 1284 -3512 1311 -3511
rect 1284 -3516 1285 -3512
rect 1289 -3516 1306 -3512
rect 1310 -3516 1311 -3512
rect 1284 -3517 1311 -3516
rect 1672 -3500 1676 -3494
rect 3076 -3446 3080 -3440
rect 3101 -3446 3106 -3390
rect 3111 -3389 3114 -3385
rect 3118 -3389 3131 -3385
rect 3135 -3389 3138 -3385
rect 3464 -3389 3468 -3379
rect 3111 -3391 3138 -3389
rect 3119 -3396 3123 -3391
rect 3127 -3446 3131 -3436
rect 3456 -3435 3460 -3429
rect 3481 -3435 3486 -3379
rect 3491 -3378 3494 -3374
rect 3498 -3378 3511 -3374
rect 3515 -3378 3518 -3374
rect 3491 -3380 3518 -3378
rect 3499 -3385 3503 -3380
rect 4231 -3420 4235 -3414
rect 4256 -3420 4261 -3364
rect 4266 -3363 4269 -3359
rect 4273 -3363 4286 -3359
rect 4290 -3363 4293 -3359
rect 4266 -3365 4293 -3363
rect 4274 -3370 4278 -3365
rect 4542 -3374 4546 -3354
rect 4569 -3374 4573 -3354
rect 4872 -3323 4876 -3318
rect 4899 -3323 4903 -3318
rect 6106 -3262 6133 -3259
rect 6106 -3266 6109 -3262
rect 6113 -3266 6126 -3262
rect 6130 -3266 6133 -3262
rect 6106 -3268 6133 -3266
rect 6114 -3273 6118 -3268
rect 8648 -3136 8675 -3133
rect 8648 -3140 8651 -3136
rect 8655 -3140 8668 -3136
rect 8672 -3140 8675 -3136
rect 8648 -3142 8675 -3140
rect 8656 -3147 8660 -3142
rect 8545 -3155 8550 -3153
rect 8510 -3160 8550 -3155
rect 8510 -3164 8516 -3163
rect 8510 -3168 8511 -3164
rect 8515 -3168 8516 -3164
rect 8510 -3171 8516 -3168
rect 8545 -3171 8550 -3160
rect 8605 -3166 8614 -3163
rect 8605 -3170 8607 -3166
rect 8611 -3170 8614 -3166
rect 8628 -3170 8641 -3167
rect 8605 -3171 8614 -3170
rect 8510 -3175 8522 -3171
rect 8510 -3185 8516 -3175
rect 8600 -3175 8614 -3171
rect 8542 -3183 8560 -3179
rect 8605 -3183 8614 -3175
rect 8510 -3189 8511 -3185
rect 8515 -3189 8516 -3185
rect 8510 -3190 8516 -3189
rect 8545 -3193 8550 -3183
rect 8605 -3187 8607 -3183
rect 8611 -3187 8614 -3183
rect 8605 -3190 8614 -3187
rect 8620 -3193 8624 -3190
rect 8574 -3197 8624 -3193
rect 8574 -3202 8578 -3197
rect 7398 -3212 7415 -3207
rect 7423 -3216 7427 -3204
rect 8510 -3207 8578 -3202
rect 8628 -3203 8632 -3190
rect 8635 -3197 8641 -3170
rect 8664 -3197 8668 -3187
rect 8635 -3202 8656 -3197
rect 8664 -3202 8675 -3197
rect 6933 -3247 6950 -3242
rect 6958 -3251 6962 -3239
rect 6537 -3256 6564 -3253
rect 6537 -3260 6540 -3256
rect 6544 -3260 6557 -3256
rect 6561 -3260 6564 -3256
rect 6537 -3262 6564 -3260
rect 6950 -3255 6962 -3251
rect 7415 -3220 7427 -3216
rect 8510 -3215 8516 -3214
rect 8510 -3219 8511 -3215
rect 8515 -3219 8516 -3215
rect 7415 -3224 7419 -3220
rect 8510 -3222 8516 -3219
rect 8545 -3222 8550 -3207
rect 8605 -3217 8614 -3214
rect 8605 -3221 8607 -3217
rect 8611 -3221 8614 -3217
rect 8605 -3222 8614 -3221
rect 6950 -3259 6954 -3255
rect 6545 -3267 6549 -3262
rect 6041 -3327 6050 -3322
rect 6073 -3323 6077 -3316
rect 6122 -3323 6126 -3313
rect 6472 -3321 6481 -3316
rect 6504 -3317 6508 -3310
rect 6553 -3317 6557 -3307
rect 6504 -3322 6545 -3317
rect 6553 -3322 6564 -3317
rect 6073 -3328 6114 -3323
rect 6122 -3328 6133 -3323
rect 6504 -3325 6508 -3322
rect 6553 -3325 6557 -3322
rect 6073 -3331 6077 -3328
rect 6122 -3331 6126 -3328
rect 6058 -3335 6095 -3331
rect 6058 -3341 6062 -3335
rect 6091 -3341 6095 -3335
rect 4588 -3373 4615 -3370
rect 4542 -3378 4583 -3374
rect 4527 -3384 4534 -3379
rect 4561 -3388 4565 -3378
rect 4282 -3420 4286 -3410
rect 4231 -3424 4245 -3420
rect 3507 -3435 3511 -3425
rect 4239 -3425 4245 -3424
rect 4256 -3425 4274 -3420
rect 4282 -3425 4295 -3420
rect 3456 -3439 3470 -3435
rect 3464 -3440 3470 -3439
rect 3481 -3440 3499 -3435
rect 3507 -3440 3520 -3435
rect 4205 -3436 4231 -3431
rect 4239 -3439 4243 -3425
rect 4282 -3428 4286 -3425
rect 3076 -3450 3090 -3446
rect 3084 -3451 3090 -3450
rect 3101 -3451 3119 -3446
rect 3127 -3451 3140 -3446
rect 3430 -3451 3456 -3446
rect 3050 -3462 3076 -3457
rect 3084 -3465 3088 -3451
rect 3127 -3454 3131 -3451
rect 3464 -3454 3468 -3440
rect 3507 -3443 3511 -3440
rect 2781 -3471 2785 -3465
rect 2773 -3472 2800 -3471
rect 2773 -3476 2774 -3472
rect 2778 -3476 2795 -3472
rect 2799 -3476 2800 -3472
rect 2773 -3477 2800 -3476
rect 1664 -3501 1691 -3500
rect 1664 -3505 1665 -3501
rect 1669 -3505 1686 -3501
rect 1690 -3505 1691 -3501
rect 2738 -3502 2742 -3496
rect 1664 -3506 1691 -3505
rect 2730 -3503 2757 -3502
rect 2730 -3507 2731 -3503
rect 2735 -3507 2752 -3503
rect 2756 -3507 2757 -3503
rect 2730 -3508 2757 -3507
rect 3119 -3480 3123 -3474
rect 3111 -3481 3138 -3480
rect 3111 -3485 3112 -3481
rect 3116 -3485 3133 -3481
rect 3137 -3485 3138 -3481
rect 3111 -3486 3138 -3485
rect 3499 -3469 3503 -3463
rect 3491 -3470 3518 -3469
rect 3491 -3474 3492 -3470
rect 3496 -3474 3513 -3470
rect 3517 -3474 3518 -3470
rect 3491 -3475 3518 -3474
rect 4553 -3434 4557 -3428
rect 4578 -3434 4583 -3378
rect 4588 -3377 4591 -3373
rect 4595 -3377 4608 -3373
rect 4612 -3377 4615 -3373
rect 4588 -3379 4615 -3377
rect 4596 -3384 4600 -3379
rect 4880 -3383 4884 -3363
rect 4907 -3383 4911 -3363
rect 5260 -3372 5264 -3352
rect 5287 -3372 5291 -3352
rect 6489 -3329 6526 -3325
rect 6489 -3335 6493 -3329
rect 6522 -3335 6526 -3329
rect 6114 -3357 6118 -3351
rect 6991 -3285 7018 -3282
rect 6991 -3289 6994 -3285
rect 6998 -3289 7011 -3285
rect 7015 -3289 7018 -3285
rect 6991 -3291 7018 -3289
rect 6999 -3296 7003 -3291
rect 8510 -3226 8522 -3222
rect 8510 -3236 8516 -3226
rect 8600 -3226 8614 -3222
rect 8542 -3234 8560 -3230
rect 8605 -3234 8614 -3226
rect 8510 -3240 8511 -3236
rect 8515 -3240 8516 -3236
rect 8510 -3241 8516 -3240
rect 7456 -3250 7483 -3247
rect 7456 -3254 7459 -3250
rect 7463 -3254 7476 -3250
rect 7480 -3254 7483 -3250
rect 7456 -3256 7483 -3254
rect 8545 -3254 8550 -3234
rect 8605 -3238 8607 -3234
rect 8611 -3238 8614 -3234
rect 8605 -3241 8614 -3238
rect 8664 -3205 8668 -3202
rect 8620 -3254 8624 -3223
rect 8656 -3231 8660 -3225
rect 8648 -3232 8675 -3231
rect 8648 -3236 8649 -3232
rect 8653 -3236 8670 -3232
rect 8674 -3236 8675 -3232
rect 8648 -3237 8675 -3236
rect 7464 -3261 7468 -3256
rect 8545 -3257 8624 -3254
rect 7391 -3315 7400 -3310
rect 7423 -3311 7427 -3304
rect 7472 -3311 7476 -3301
rect 7423 -3316 7464 -3311
rect 7472 -3316 7483 -3311
rect 7423 -3319 7427 -3316
rect 7472 -3319 7476 -3316
rect 7408 -3323 7445 -3319
rect 7408 -3329 7412 -3323
rect 7441 -3329 7445 -3323
rect 6545 -3351 6549 -3345
rect 6926 -3350 6935 -3345
rect 6958 -3346 6962 -3339
rect 7007 -3346 7011 -3336
rect 6958 -3351 6999 -3346
rect 7007 -3351 7018 -3346
rect 7464 -3345 7468 -3339
rect 7456 -3346 7483 -3345
rect 6537 -3352 6564 -3351
rect 6106 -3358 6133 -3357
rect 6050 -3367 6054 -3361
rect 6083 -3367 6087 -3361
rect 6106 -3362 6107 -3358
rect 6111 -3362 6128 -3358
rect 6132 -3362 6133 -3358
rect 6481 -3361 6485 -3355
rect 6514 -3361 6518 -3355
rect 6537 -3356 6538 -3352
rect 6542 -3356 6559 -3352
rect 6563 -3356 6564 -3352
rect 6958 -3354 6962 -3351
rect 7007 -3354 7011 -3351
rect 6537 -3357 6564 -3356
rect 6943 -3358 6980 -3354
rect 6106 -3363 6133 -3362
rect 6473 -3362 6500 -3361
rect 6473 -3366 6474 -3362
rect 6478 -3366 6495 -3362
rect 6499 -3366 6500 -3362
rect 6473 -3367 6500 -3366
rect 6506 -3362 6533 -3361
rect 6506 -3366 6507 -3362
rect 6511 -3366 6528 -3362
rect 6532 -3366 6533 -3362
rect 6943 -3364 6947 -3358
rect 6976 -3364 6980 -3358
rect 6506 -3367 6533 -3366
rect 6042 -3368 6069 -3367
rect 5306 -3371 5333 -3368
rect 5260 -3376 5301 -3372
rect 4926 -3382 4953 -3379
rect 5245 -3382 5252 -3377
rect 4880 -3387 4921 -3383
rect 4865 -3393 4872 -3388
rect 4899 -3397 4903 -3387
rect 4604 -3434 4608 -3424
rect 4553 -3438 4567 -3434
rect 4561 -3439 4567 -3438
rect 4578 -3439 4596 -3434
rect 4604 -3439 4617 -3434
rect 4274 -3454 4278 -3448
rect 4527 -3450 4553 -3445
rect 4561 -3453 4565 -3439
rect 4604 -3442 4608 -3439
rect 4266 -3455 4293 -3454
rect 4266 -3459 4267 -3455
rect 4271 -3459 4288 -3455
rect 4292 -3459 4293 -3455
rect 4266 -3460 4293 -3459
rect 4231 -3485 4235 -3479
rect 4223 -3486 4250 -3485
rect 4223 -3490 4224 -3486
rect 4228 -3490 4245 -3486
rect 4249 -3490 4250 -3486
rect 4223 -3491 4250 -3490
rect 4891 -3443 4895 -3437
rect 4916 -3443 4921 -3387
rect 4926 -3386 4929 -3382
rect 4933 -3386 4946 -3382
rect 4950 -3386 4953 -3382
rect 5279 -3386 5283 -3376
rect 4926 -3388 4953 -3386
rect 4934 -3393 4938 -3388
rect 4942 -3443 4946 -3433
rect 5271 -3432 5275 -3426
rect 5296 -3432 5301 -3376
rect 5306 -3375 5309 -3371
rect 5313 -3375 5326 -3371
rect 5330 -3375 5333 -3371
rect 6042 -3372 6043 -3368
rect 6047 -3372 6064 -3368
rect 6068 -3372 6069 -3368
rect 6042 -3373 6069 -3372
rect 6075 -3368 6102 -3367
rect 6075 -3372 6076 -3368
rect 6080 -3372 6097 -3368
rect 6101 -3372 6102 -3368
rect 6075 -3373 6102 -3372
rect 5306 -3377 5333 -3375
rect 5314 -3382 5318 -3377
rect 7400 -3355 7404 -3349
rect 7433 -3355 7437 -3349
rect 7456 -3350 7457 -3346
rect 7461 -3350 7478 -3346
rect 7482 -3350 7483 -3346
rect 7456 -3351 7483 -3350
rect 7392 -3356 7419 -3355
rect 7392 -3360 7393 -3356
rect 7397 -3360 7414 -3356
rect 7418 -3360 7419 -3356
rect 7392 -3361 7419 -3360
rect 7425 -3356 7452 -3355
rect 7425 -3360 7426 -3356
rect 7430 -3360 7447 -3356
rect 7451 -3360 7452 -3356
rect 7425 -3361 7452 -3360
rect 6999 -3380 7003 -3374
rect 6991 -3381 7018 -3380
rect 6935 -3390 6939 -3384
rect 6968 -3390 6972 -3384
rect 6991 -3385 6992 -3381
rect 6996 -3385 7013 -3381
rect 7017 -3385 7018 -3381
rect 6991 -3386 7018 -3385
rect 6927 -3391 6954 -3390
rect 6927 -3395 6928 -3391
rect 6932 -3395 6949 -3391
rect 6953 -3395 6954 -3391
rect 6927 -3396 6954 -3395
rect 6960 -3391 6987 -3390
rect 6960 -3395 6961 -3391
rect 6965 -3395 6982 -3391
rect 6986 -3395 6987 -3391
rect 6960 -3396 6987 -3395
rect 5322 -3432 5326 -3422
rect 5271 -3436 5285 -3432
rect 5279 -3437 5285 -3436
rect 5296 -3437 5314 -3432
rect 5322 -3437 5335 -3432
rect 4891 -3447 4905 -3443
rect 4899 -3448 4905 -3447
rect 4916 -3448 4934 -3443
rect 4942 -3448 4955 -3443
rect 5245 -3448 5271 -3443
rect 4865 -3459 4891 -3454
rect 4899 -3462 4903 -3448
rect 4942 -3451 4946 -3448
rect 5279 -3451 5283 -3437
rect 5322 -3440 5326 -3437
rect 4596 -3468 4600 -3462
rect 4588 -3469 4615 -3468
rect 4588 -3473 4589 -3469
rect 4593 -3473 4610 -3469
rect 4614 -3473 4615 -3469
rect 4588 -3474 4615 -3473
rect 3456 -3500 3460 -3494
rect 4553 -3499 4557 -3493
rect 4545 -3500 4572 -3499
rect 3448 -3501 3475 -3500
rect 3448 -3505 3449 -3501
rect 3453 -3505 3470 -3501
rect 3474 -3505 3475 -3501
rect 4545 -3504 4546 -3500
rect 4550 -3504 4567 -3500
rect 4571 -3504 4572 -3500
rect 4545 -3505 4572 -3504
rect 4934 -3477 4938 -3471
rect 4926 -3478 4953 -3477
rect 4926 -3482 4927 -3478
rect 4931 -3482 4948 -3478
rect 4952 -3482 4953 -3478
rect 4926 -3483 4953 -3482
rect 5314 -3466 5318 -3460
rect 5306 -3467 5333 -3466
rect 5306 -3471 5307 -3467
rect 5311 -3471 5328 -3467
rect 5332 -3471 5333 -3467
rect 5306 -3472 5333 -3471
rect 5271 -3497 5275 -3491
rect 5263 -3498 5290 -3497
rect 5263 -3502 5264 -3498
rect 5268 -3502 5285 -3498
rect 5289 -3502 5290 -3498
rect 3076 -3511 3080 -3505
rect 3448 -3506 3475 -3505
rect 4891 -3508 4895 -3502
rect 5263 -3503 5290 -3502
rect 4883 -3509 4910 -3508
rect 3068 -3512 3095 -3511
rect 3068 -3516 3069 -3512
rect 3073 -3516 3090 -3512
rect 3094 -3516 3095 -3512
rect 4883 -3513 4884 -3509
rect 4888 -3513 4905 -3509
rect 4909 -3513 4910 -3509
rect 4883 -3514 4910 -3513
rect 3068 -3517 3095 -3516
rect 1629 -3531 1633 -3525
rect 1621 -3532 1648 -3531
rect 1621 -3536 1622 -3532
rect 1626 -3536 1643 -3532
rect 1647 -3536 1648 -3532
rect 1249 -3542 1253 -3536
rect 1621 -3537 1648 -3536
rect 1241 -3543 1268 -3542
rect 1241 -3547 1242 -3543
rect 1246 -3547 1263 -3543
rect 1267 -3547 1268 -3543
rect 1241 -3548 1268 -3547
rect 59 -3583 63 -3563
rect 86 -3583 90 -3563
rect 105 -3582 132 -3579
rect 59 -3587 100 -3583
rect -27 -3593 51 -3588
rect -27 -3594 -18 -3593
rect 78 -3597 82 -3587
rect 70 -3643 74 -3637
rect 95 -3643 100 -3587
rect 105 -3586 108 -3582
rect 112 -3586 125 -3582
rect 129 -3586 132 -3582
rect 105 -3588 132 -3586
rect 113 -3593 117 -3588
rect 121 -3643 125 -3633
rect 70 -3647 84 -3643
rect 78 -3648 84 -3647
rect 95 -3648 113 -3643
rect 121 -3648 134 -3643
rect -52 -3659 70 -3654
rect 78 -3662 82 -3648
rect 121 -3651 125 -3648
rect 113 -3677 117 -3671
rect 105 -3678 132 -3677
rect 105 -3682 106 -3678
rect 110 -3682 127 -3678
rect 131 -3682 132 -3678
rect 105 -3683 132 -3682
rect 70 -3708 74 -3702
rect 62 -3709 89 -3708
rect 62 -3713 63 -3709
rect 67 -3713 84 -3709
rect 88 -3713 89 -3709
rect 62 -3714 89 -3713
<< m2contact >>
rect -842 514 -833 519
rect -32 -75 -23 -70
rect -12 -868 -3 -863
rect -27 -1992 -18 -1987
rect -27 -3411 -18 -3406
<< metal2 >>
rect -917 514 -842 519
rect -107 -75 -32 -70
rect -87 -868 -12 -863
rect -102 -1992 -27 -1987
rect -102 -3411 -27 -3406
<< labels >>
rlabel metal1 -61 254 -61 254 7 vdd
rlabel metal1 -157 254 -157 254 3 gnd
rlabel metal1 -61 305 -61 305 7 vdd
rlabel metal1 -157 305 -157 305 3 gnd
rlabel metal1 -9 247 -9 247 1 gnd
rlabel metal1 -9 343 -9 343 5 vdd
rlabel metal1 318 192 318 192 1 gnd
rlabel metal1 318 288 318 288 5 vdd
rlabel metal1 275 161 275 161 1 gnd
rlabel metal1 283 358 283 358 5 vdd
rlabel metal1 256 358 256 358 5 vdd
rlabel metal1 82 231 82 231 1 gnd
rlabel metal1 82 327 82 327 5 vdd
rlabel metal1 691 -382 691 -382 1 gnd
rlabel metal1 691 -286 691 -286 5 vdd
rlabel metal1 648 -413 648 -413 1 gnd
rlabel metal1 656 -216 656 -216 5 vdd
rlabel metal1 629 -216 629 -216 5 vdd
rlabel metal1 147 370 147 370 5 vdd
rlabel metal1 132 127 132 127 1 gnd
rlabel metal1 165 127 165 127 1 gnd
rlabel metal1 196 233 196 233 5 vdd
rlabel metal1 196 137 196 137 1 gnd
rlabel metal1 926 -158 926 -158 5 vdd
rlabel metal1 911 -401 911 -401 1 gnd
rlabel metal1 944 -401 944 -401 1 gnd
rlabel metal1 975 -295 975 -295 5 vdd
rlabel metal1 975 -391 975 -391 1 gnd
rlabel metal1 1329 -40 1329 -40 7 vdd
rlabel metal1 1233 -40 1233 -40 3 gnd
rlabel metal1 1329 11 1329 11 7 vdd
rlabel metal1 1233 11 1233 11 3 gnd
rlabel metal1 1381 -47 1381 -47 1 gnd
rlabel metal1 1381 49 1381 49 5 vdd
rlabel metal1 122 -888 122 -888 7 vdd
rlabel metal1 26 -888 26 -888 3 gnd
rlabel metal1 122 -837 122 -837 7 vdd
rlabel metal1 26 -837 26 -837 3 gnd
rlabel metal1 174 -895 174 -895 1 gnd
rlabel metal1 174 -799 174 -799 5 vdd
rlabel metal1 133 -1137 133 -1137 1 gnd
rlabel metal1 133 -1041 133 -1041 5 vdd
rlabel metal1 90 -1168 90 -1168 1 gnd
rlabel metal1 98 -971 98 -971 5 vdd
rlabel metal1 71 -971 71 -971 5 vdd
rlabel metal1 -708 494 -708 494 7 vdd
rlabel metal1 -804 494 -804 494 3 gnd
rlabel metal1 -708 545 -708 545 7 vdd
rlabel metal1 -804 545 -804 545 3 gnd
rlabel metal1 -656 487 -656 487 1 gnd
rlabel metal1 -656 583 -656 583 5 vdd
rlabel metal1 -697 245 -697 245 1 gnd
rlabel metal1 -697 341 -697 341 5 vdd
rlabel metal1 -740 214 -740 214 1 gnd
rlabel metal1 -732 411 -732 411 5 vdd
rlabel metal1 -759 411 -759 411 5 vdd
rlabel metal1 102 -95 102 -95 7 vdd
rlabel metal1 6 -95 6 -95 3 gnd
rlabel metal1 102 -44 102 -44 7 vdd
rlabel metal1 6 -44 6 -44 3 gnd
rlabel metal1 154 -102 154 -102 1 gnd
rlabel metal1 154 -6 154 -6 5 vdd
rlabel metal1 113 -344 113 -344 1 gnd
rlabel metal1 113 -248 113 -248 5 vdd
rlabel metal1 70 -375 70 -375 1 gnd
rlabel metal1 78 -178 78 -178 5 vdd
rlabel metal1 51 -178 51 -178 5 vdd
rlabel metal1 56 -2095 56 -2095 5 vdd
rlabel metal1 83 -2095 83 -2095 5 vdd
rlabel metal1 75 -2292 75 -2292 1 gnd
rlabel metal1 118 -2165 118 -2165 5 vdd
rlabel metal1 118 -2261 118 -2261 1 gnd
rlabel metal1 159 -1923 159 -1923 5 vdd
rlabel metal1 159 -2019 159 -2019 1 gnd
rlabel metal1 11 -1961 11 -1961 3 gnd
rlabel metal1 107 -1961 107 -1961 7 vdd
rlabel metal1 11 -2012 11 -2012 3 gnd
rlabel metal1 107 -2012 107 -2012 7 vdd
rlabel metal1 56 -3514 56 -3514 5 vdd
rlabel metal1 83 -3514 83 -3514 5 vdd
rlabel metal1 75 -3711 75 -3711 1 gnd
rlabel metal1 118 -3584 118 -3584 5 vdd
rlabel metal1 118 -3680 118 -3680 1 gnd
rlabel metal1 159 -3342 159 -3342 5 vdd
rlabel metal1 159 -3438 159 -3438 1 gnd
rlabel metal1 11 -3380 11 -3380 3 gnd
rlabel metal1 107 -3380 107 -3380 7 vdd
rlabel metal1 11 -3431 11 -3431 3 gnd
rlabel metal1 107 -3431 107 -3431 7 vdd
rlabel metal1 734 -1018 734 -1018 1 gnd
rlabel metal1 734 -922 734 -922 5 vdd
rlabel metal1 691 -1049 691 -1049 1 gnd
rlabel metal1 699 -852 699 -852 5 vdd
rlabel metal1 672 -852 672 -852 5 vdd
rlabel metal1 1072 -1027 1072 -1027 1 gnd
rlabel metal1 1072 -931 1072 -931 5 vdd
rlabel metal1 1029 -1058 1029 -1058 1 gnd
rlabel metal1 1037 -861 1037 -861 5 vdd
rlabel metal1 1010 -861 1010 -861 5 vdd
rlabel metal1 1390 -850 1390 -850 5 vdd
rlabel metal1 1417 -850 1417 -850 5 vdd
rlabel metal1 1409 -1047 1409 -1047 1 gnd
rlabel metal1 1452 -920 1452 -920 5 vdd
rlabel metal1 1452 -1016 1452 -1016 1 gnd
rlabel metal1 806 -1913 806 -1913 5 vdd
rlabel metal1 833 -1913 833 -1913 5 vdd
rlabel metal1 825 -2110 825 -2110 1 gnd
rlabel metal1 868 -1983 868 -1983 5 vdd
rlabel metal1 868 -2079 868 -2079 1 gnd
rlabel metal1 1274 -1904 1274 -1904 5 vdd
rlabel metal1 1301 -1904 1301 -1904 5 vdd
rlabel metal1 1293 -2101 1293 -2101 1 gnd
rlabel metal1 1336 -1974 1336 -1974 5 vdd
rlabel metal1 1336 -2070 1336 -2070 1 gnd
rlabel metal1 1676 -1901 1676 -1901 5 vdd
rlabel metal1 1703 -1901 1703 -1901 5 vdd
rlabel metal1 1695 -2098 1695 -2098 1 gnd
rlabel metal1 1738 -1971 1738 -1971 5 vdd
rlabel metal1 1738 -2067 1738 -2067 1 gnd
rlabel metal1 2177 -1866 2177 -1866 5 vdd
rlabel metal1 2204 -1866 2204 -1866 5 vdd
rlabel metal1 2196 -2063 2196 -2063 1 gnd
rlabel metal1 2239 -1936 2239 -1936 5 vdd
rlabel metal1 2239 -2032 2239 -2032 1 gnd
rlabel metal1 2782 -1866 2782 -1866 5 vdd
rlabel metal1 2809 -1866 2809 -1866 5 vdd
rlabel metal1 2801 -2063 2801 -2063 1 gnd
rlabel metal1 2844 -1936 2844 -1936 5 vdd
rlabel metal1 2844 -2032 2844 -2032 1 gnd
rlabel metal1 3387 -1866 3387 -1866 5 vdd
rlabel metal1 3414 -1866 3414 -1866 5 vdd
rlabel metal1 3406 -2063 3406 -2063 1 gnd
rlabel metal1 3449 -1936 3449 -1936 5 vdd
rlabel metal1 3449 -2032 3449 -2032 1 gnd
rlabel metal1 959 -3505 959 -3505 1 gnd
rlabel metal1 959 -3409 959 -3409 5 vdd
rlabel metal1 916 -3536 916 -3536 1 gnd
rlabel metal1 924 -3339 924 -3339 5 vdd
rlabel metal1 897 -3339 897 -3339 5 vdd
rlabel metal1 1297 -3514 1297 -3514 1 gnd
rlabel metal1 1297 -3418 1297 -3418 5 vdd
rlabel metal1 1254 -3545 1254 -3545 1 gnd
rlabel metal1 1262 -3348 1262 -3348 5 vdd
rlabel metal1 1235 -3348 1235 -3348 5 vdd
rlabel metal1 1615 -3337 1615 -3337 5 vdd
rlabel metal1 1642 -3337 1642 -3337 5 vdd
rlabel metal1 1634 -3534 1634 -3534 1 gnd
rlabel metal1 1677 -3407 1677 -3407 5 vdd
rlabel metal1 1677 -3503 1677 -3503 1 gnd
rlabel metal1 2786 -3474 2786 -3474 1 gnd
rlabel metal1 2786 -3378 2786 -3378 5 vdd
rlabel metal1 2743 -3505 2743 -3505 1 gnd
rlabel metal1 2751 -3308 2751 -3308 5 vdd
rlabel metal1 2724 -3308 2724 -3308 5 vdd
rlabel metal1 3124 -3483 3124 -3483 1 gnd
rlabel metal1 3124 -3387 3124 -3387 5 vdd
rlabel metal1 3081 -3514 3081 -3514 1 gnd
rlabel metal1 3089 -3317 3089 -3317 5 vdd
rlabel metal1 3062 -3317 3062 -3317 5 vdd
rlabel metal1 3442 -3306 3442 -3306 5 vdd
rlabel metal1 3469 -3306 3469 -3306 5 vdd
rlabel metal1 3461 -3503 3461 -3503 1 gnd
rlabel metal1 3504 -3376 3504 -3376 5 vdd
rlabel metal1 3504 -3472 3504 -3472 1 gnd
rlabel metal1 4601 -3471 4601 -3471 1 gnd
rlabel metal1 4601 -3375 4601 -3375 5 vdd
rlabel metal1 4558 -3502 4558 -3502 1 gnd
rlabel metal1 4566 -3305 4566 -3305 5 vdd
rlabel metal1 4539 -3305 4539 -3305 5 vdd
rlabel metal1 4939 -3480 4939 -3480 1 gnd
rlabel metal1 4939 -3384 4939 -3384 5 vdd
rlabel metal1 4896 -3511 4896 -3511 1 gnd
rlabel metal1 4904 -3314 4904 -3314 5 vdd
rlabel metal1 4877 -3314 4877 -3314 5 vdd
rlabel metal1 5257 -3303 5257 -3303 5 vdd
rlabel metal1 5284 -3303 5284 -3303 5 vdd
rlabel metal1 5276 -3500 5276 -3500 1 gnd
rlabel metal1 5319 -3373 5319 -3373 5 vdd
rlabel metal1 5319 -3469 5319 -3469 1 gnd
rlabel metal1 4279 -3457 4279 -3457 1 gnd
rlabel metal1 4279 -3361 4279 -3361 5 vdd
rlabel metal1 4236 -3488 4236 -3488 1 gnd
rlabel metal1 4244 -3291 4244 -3291 5 vdd
rlabel metal1 4217 -3291 4217 -3291 5 vdd
rlabel metal1 2232 -663 2232 -663 5 vdd
rlabel metal1 2217 -906 2217 -906 1 gnd
rlabel metal1 2250 -906 2250 -906 1 gnd
rlabel metal1 2281 -800 2281 -800 5 vdd
rlabel metal1 2281 -896 2281 -896 1 gnd
rlabel metal1 2726 -646 2726 -646 5 vdd
rlabel metal1 2711 -889 2711 -889 1 gnd
rlabel metal1 2744 -889 2744 -889 1 gnd
rlabel metal1 2775 -783 2775 -783 5 vdd
rlabel metal1 2775 -879 2775 -879 1 gnd
rlabel metal1 4064 -2003 4064 -2003 1 gnd
rlabel metal1 4064 -1907 4064 -1907 5 vdd
rlabel metal1 4033 -2013 4033 -2013 1 gnd
rlabel metal1 4000 -2013 4000 -2013 1 gnd
rlabel metal1 4015 -1770 4015 -1770 5 vdd
rlabel metal1 4518 -2032 4518 -2032 1 gnd
rlabel metal1 4518 -1936 4518 -1936 5 vdd
rlabel metal1 4487 -2042 4487 -2042 1 gnd
rlabel metal1 4454 -2042 4454 -2042 1 gnd
rlabel metal1 4469 -1799 4469 -1799 5 vdd
rlabel metal1 4983 -1997 4983 -1997 1 gnd
rlabel metal1 4983 -1901 4983 -1901 5 vdd
rlabel metal1 4952 -2007 4952 -2007 1 gnd
rlabel metal1 4919 -2007 4919 -2007 1 gnd
rlabel metal1 4934 -1764 4934 -1764 5 vdd
rlabel metal1 6119 -3360 6119 -3360 1 gnd
rlabel metal1 6119 -3264 6119 -3264 5 vdd
rlabel metal1 6088 -3370 6088 -3370 1 gnd
rlabel metal1 6055 -3370 6055 -3370 1 gnd
rlabel metal1 6070 -3127 6070 -3127 5 vdd
rlabel metal1 6550 -3354 6550 -3354 1 gnd
rlabel metal1 6550 -3258 6550 -3258 5 vdd
rlabel metal1 6519 -3364 6519 -3364 1 gnd
rlabel metal1 6486 -3364 6486 -3364 1 gnd
rlabel metal1 6501 -3121 6501 -3121 5 vdd
rlabel metal1 7004 -3383 7004 -3383 1 gnd
rlabel metal1 7004 -3287 7004 -3287 5 vdd
rlabel metal1 6973 -3393 6973 -3393 1 gnd
rlabel metal1 6940 -3393 6940 -3393 1 gnd
rlabel metal1 6955 -3150 6955 -3150 5 vdd
rlabel metal1 7469 -3348 7469 -3348 1 gnd
rlabel metal1 7469 -3252 7469 -3252 5 vdd
rlabel metal1 7438 -3358 7438 -3358 1 gnd
rlabel metal1 7405 -3358 7405 -3358 1 gnd
rlabel metal1 7420 -3115 7420 -3115 5 vdd
rlabel metal1 3661 -628 3661 -628 5 vdd
rlabel metal1 3661 -724 3661 -724 1 gnd
rlabel metal1 3513 -666 3513 -666 3 gnd
rlabel metal1 3609 -666 3609 -666 7 vdd
rlabel metal1 3513 -717 3513 -717 3 gnd
rlabel metal1 3609 -717 3609 -717 7 vdd
rlabel metal1 5987 -1723 5987 -1723 5 vdd
rlabel metal1 5987 -1819 5987 -1819 1 gnd
rlabel metal1 5839 -1761 5839 -1761 3 gnd
rlabel metal1 5935 -1761 5935 -1761 7 vdd
rlabel metal1 5839 -1812 5839 -1812 3 gnd
rlabel metal1 5935 -1812 5935 -1812 7 vdd
rlabel metal1 8661 -3138 8661 -3138 5 vdd
rlabel metal1 8661 -3234 8661 -3234 1 gnd
rlabel metal1 8513 -3176 8513 -3176 3 gnd
rlabel metal1 8609 -3176 8609 -3176 7 vdd
rlabel metal1 8513 -3227 8513 -3227 3 gnd
rlabel metal1 8609 -3227 8609 -3227 7 vdd
<< end >>
