magic
tech scmos
timestamp 1731863020
<< nwell >>
rect 804 1631 866 1658
rect 900 1626 927 1688
rect 991 1610 1018 1672
rect 804 1580 866 1607
rect 1056 1513 1083 1715
rect 1165 1641 1219 1703
rect 1105 1516 1132 1578
rect 1227 1571 1254 1633
rect 2852 1604 2914 1631
rect 2948 1599 2975 1661
rect 3039 1583 3066 1645
rect 2852 1553 2914 1580
rect 3104 1486 3131 1688
rect 3213 1614 3267 1676
rect 3153 1489 3180 1551
rect 3275 1544 3302 1606
rect -1538 288 -1506 414
rect -1486 288 -1454 414
rect -1434 350 -1402 414
rect -1382 350 -1350 414
rect -1337 358 -1273 422
rect 3757 285 3789 411
rect 3809 285 3841 411
rect 3861 347 3893 411
rect 3913 347 3945 411
rect 3958 355 4022 419
rect -412 -113 -380 13
rect -360 -113 -328 13
rect -308 -51 -276 13
rect -256 -51 -224 13
rect -211 -43 -147 21
rect 1063 -7 1125 20
rect 1159 -12 1186 50
rect 1409 -18 1441 108
rect 1461 -18 1493 108
rect 1513 44 1545 108
rect 1565 44 1597 108
rect 1610 52 1674 116
rect 150 -206 212 -179
rect 246 -211 273 -149
rect 438 -193 492 -131
rect -416 -368 -384 -242
rect -364 -368 -332 -242
rect -312 -306 -280 -242
rect -260 -306 -228 -242
rect -215 -298 -151 -234
rect 150 -257 212 -230
rect 500 -263 527 -201
rect 808 -248 835 -46
rect 1063 -58 1125 -31
rect 857 -245 884 -183
rect 1058 -227 1120 -200
rect 1154 -232 1181 -170
rect 1058 -278 1120 -251
rect 163 -355 217 -293
rect 1424 -294 1456 -168
rect 1476 -294 1508 -168
rect 1528 -232 1560 -168
rect 1580 -232 1612 -168
rect 1625 -224 1689 -160
rect 225 -425 252 -363
rect -319 -950 -287 -824
rect -267 -950 -235 -824
rect -215 -888 -183 -824
rect -163 -888 -131 -824
rect -118 -880 -54 -816
rect 618 -844 672 -782
rect 680 -914 707 -852
rect 952 -895 979 -693
rect 1001 -892 1028 -830
rect 1203 -897 1230 -695
rect 1252 -894 1279 -832
rect 138 -992 200 -965
rect 234 -997 261 -935
rect 1510 -957 1572 -930
rect 1606 -962 1633 -900
rect 1808 -967 1840 -841
rect 1860 -967 1892 -841
rect 1912 -905 1944 -841
rect 1964 -905 1996 -841
rect 2009 -897 2073 -833
rect 1510 -1008 1572 -981
rect -3549 -1226 -3487 -1199
rect -3453 -1231 -3426 -1169
rect -3362 -1247 -3335 -1185
rect -3549 -1277 -3487 -1250
rect -3297 -1344 -3270 -1142
rect -3188 -1216 -3134 -1154
rect -338 -1173 -306 -1047
rect -286 -1173 -254 -1047
rect -234 -1111 -202 -1047
rect -182 -1111 -150 -1047
rect -137 -1103 -73 -1039
rect 138 -1043 200 -1016
rect 151 -1141 205 -1079
rect 541 -1089 595 -1027
rect 759 -1089 813 -1027
rect 213 -1211 240 -1149
rect 603 -1159 630 -1097
rect 821 -1159 848 -1097
rect -3248 -1341 -3221 -1279
rect -3126 -1286 -3099 -1224
rect -338 -1511 -306 -1385
rect -286 -1511 -254 -1385
rect -234 -1449 -202 -1385
rect -182 -1449 -150 -1385
rect -137 -1441 -73 -1377
rect 553 -1404 607 -1342
rect 615 -1474 642 -1412
rect 147 -1652 209 -1625
rect 243 -1657 270 -1595
rect 147 -1703 209 -1676
rect 554 -1687 608 -1625
rect 790 -1634 844 -1572
rect 1072 -1620 1099 -1418
rect 1121 -1617 1148 -1555
rect -353 -1848 -321 -1722
rect -301 -1848 -269 -1722
rect -249 -1786 -217 -1722
rect -197 -1786 -165 -1722
rect -152 -1778 -88 -1714
rect 160 -1801 214 -1739
rect 616 -1757 643 -1695
rect 852 -1704 879 -1642
rect 222 -1871 249 -1809
rect 799 -1845 853 -1783
rect 550 -1958 604 -1896
rect 861 -1915 888 -1853
rect 1083 -1920 1110 -1718
rect 1369 -1773 1396 -1571
rect 1691 -1693 1753 -1666
rect 1787 -1698 1814 -1636
rect 1418 -1770 1445 -1708
rect 1997 -1717 2029 -1591
rect 2049 -1717 2081 -1591
rect 2101 -1655 2133 -1591
rect 2153 -1655 2185 -1591
rect 2198 -1647 2262 -1583
rect 1691 -1744 1753 -1717
rect 1132 -1917 1159 -1855
rect 612 -2028 639 -1966
rect 538 -2207 592 -2145
rect 600 -2277 627 -2215
rect -353 -2455 -321 -2329
rect -301 -2455 -269 -2329
rect -249 -2393 -217 -2329
rect -197 -2393 -165 -2329
rect -152 -2385 -88 -2321
rect 144 -2527 206 -2500
rect 240 -2532 267 -2470
rect 144 -2578 206 -2551
rect 631 -2554 685 -2492
rect -353 -2725 -321 -2599
rect -301 -2725 -269 -2599
rect -249 -2663 -217 -2599
rect -197 -2663 -165 -2599
rect -152 -2655 -88 -2591
rect 157 -2676 211 -2614
rect 693 -2624 720 -2562
rect 966 -2606 1020 -2544
rect 1028 -2676 1055 -2614
rect 219 -2746 246 -2684
rect 1296 -2687 1323 -2485
rect 1345 -2684 1372 -2622
rect 632 -2837 686 -2775
rect 694 -2907 721 -2845
rect 967 -2889 1021 -2827
rect 1029 -2959 1056 -2897
rect 628 -3108 682 -3046
rect 1303 -3076 1330 -2874
rect 1800 -3001 1827 -2799
rect 1849 -2998 1876 -2936
rect 2071 -2959 2103 -2833
rect 2123 -2959 2155 -2833
rect 2175 -2897 2207 -2833
rect 2227 -2897 2259 -2833
rect 2272 -2889 2336 -2825
rect 1352 -3073 1379 -3011
rect 690 -3178 717 -3116
rect 1297 -3291 1351 -3229
rect 1595 -3232 1622 -3030
rect 1644 -3229 1671 -3167
rect 616 -3357 670 -3295
rect 1359 -3361 1386 -3299
rect 678 -3427 705 -3365
rect 957 -3423 1011 -3361
rect 1019 -3493 1046 -3431
rect 633 -3624 687 -3562
rect 695 -3694 722 -3632
rect 621 -3873 675 -3811
rect 683 -3943 710 -3881
<< ntransistor >>
rect 774 1643 794 1645
rect 877 1631 879 1651
rect 877 1598 879 1618
rect 913 1596 915 1616
rect 774 1592 794 1594
rect 1004 1580 1006 1600
rect 1197 1575 1199 1615
rect 2822 1616 2842 1618
rect 2925 1604 2927 1624
rect 2925 1571 2927 1591
rect 2961 1569 2963 1589
rect 2822 1565 2842 1567
rect 1197 1510 1199 1550
rect 1240 1541 1242 1561
rect 3052 1553 3054 1573
rect 1054 1476 1056 1496
rect 1087 1476 1089 1496
rect 1118 1486 1120 1506
rect 3245 1548 3247 1588
rect 3245 1483 3247 1523
rect 3288 1514 3290 1534
rect 3102 1449 3104 1469
rect 3135 1449 3137 1469
rect 3166 1459 3168 1479
rect -1322 327 -1320 347
rect -1290 327 -1288 347
rect -1419 303 -1417 323
rect -1367 303 -1365 323
rect 3973 324 3975 344
rect 4005 324 4007 344
rect 3876 300 3878 320
rect 3928 300 3930 320
rect -1523 256 -1521 276
rect -1471 256 -1469 276
rect -1419 256 -1417 276
rect -1367 256 -1365 276
rect 3772 253 3774 273
rect 3824 253 3826 273
rect 3876 253 3878 273
rect 3928 253 3930 273
rect 1033 5 1053 7
rect 1136 -7 1138 13
rect 1136 -40 1138 -20
rect 1625 21 1627 41
rect 1657 21 1659 41
rect 1528 -3 1530 17
rect 1580 -3 1582 17
rect 1172 -42 1174 -22
rect 1033 -46 1053 -44
rect -196 -74 -194 -54
rect -164 -74 -162 -54
rect 1424 -50 1426 -30
rect 1476 -50 1478 -30
rect 1528 -50 1530 -30
rect 1580 -50 1582 -30
rect -293 -98 -291 -78
rect -241 -98 -239 -78
rect -397 -145 -395 -125
rect -345 -145 -343 -125
rect -293 -145 -291 -125
rect -241 -145 -239 -125
rect 120 -194 140 -192
rect 223 -206 225 -186
rect 223 -239 225 -219
rect 259 -241 261 -221
rect 120 -245 140 -243
rect 470 -259 472 -219
rect 1028 -215 1048 -213
rect 1131 -227 1133 -207
rect -200 -329 -198 -309
rect -168 -329 -166 -309
rect -297 -353 -295 -333
rect -245 -353 -243 -333
rect 470 -324 472 -284
rect 513 -293 515 -273
rect 806 -285 808 -265
rect 839 -285 841 -265
rect 870 -275 872 -255
rect 1131 -260 1133 -240
rect 1167 -262 1169 -242
rect 1028 -266 1048 -264
rect 1640 -255 1642 -235
rect 1672 -255 1674 -235
rect 1543 -279 1545 -259
rect 1595 -279 1597 -259
rect 1439 -326 1441 -306
rect 1491 -326 1493 -306
rect 1543 -326 1545 -306
rect 1595 -326 1597 -306
rect -401 -400 -399 -380
rect -349 -400 -347 -380
rect -297 -400 -295 -380
rect -245 -400 -243 -380
rect 195 -421 197 -381
rect 195 -486 197 -446
rect 238 -455 240 -435
rect -103 -911 -101 -891
rect -71 -911 -69 -891
rect 650 -910 652 -870
rect -200 -935 -198 -915
rect -148 -935 -146 -915
rect -304 -982 -302 -962
rect -252 -982 -250 -962
rect -200 -982 -198 -962
rect -148 -982 -146 -962
rect 108 -980 128 -978
rect 211 -992 213 -972
rect 650 -975 652 -935
rect 693 -944 695 -924
rect 950 -932 952 -912
rect 983 -932 985 -912
rect 1014 -922 1016 -902
rect 1201 -934 1203 -914
rect 1234 -934 1236 -914
rect 1265 -924 1267 -904
rect 1480 -945 1500 -943
rect 1583 -957 1585 -937
rect 211 -1025 213 -1005
rect 1583 -990 1585 -970
rect 2024 -928 2026 -908
rect 2056 -928 2058 -908
rect 1927 -952 1929 -932
rect 1979 -952 1981 -932
rect 1619 -992 1621 -972
rect 1480 -996 1500 -994
rect 1823 -999 1825 -979
rect 1875 -999 1877 -979
rect 1927 -999 1929 -979
rect 1979 -999 1981 -979
rect 247 -1027 249 -1007
rect 108 -1031 128 -1029
rect -3579 -1214 -3559 -1212
rect -3476 -1226 -3474 -1206
rect -3476 -1259 -3474 -1239
rect -122 -1134 -120 -1114
rect -90 -1134 -88 -1114
rect -219 -1158 -217 -1138
rect -167 -1158 -165 -1138
rect -323 -1205 -321 -1185
rect -271 -1205 -269 -1185
rect -219 -1205 -217 -1185
rect -167 -1205 -165 -1185
rect -3440 -1261 -3438 -1241
rect 183 -1207 185 -1167
rect -3579 -1265 -3559 -1263
rect -3349 -1277 -3347 -1257
rect -3156 -1282 -3154 -1242
rect 573 -1155 575 -1115
rect 791 -1155 793 -1115
rect 573 -1220 575 -1180
rect 616 -1189 618 -1169
rect 791 -1220 793 -1180
rect 834 -1189 836 -1169
rect 183 -1272 185 -1232
rect 226 -1241 228 -1221
rect -3156 -1347 -3154 -1307
rect -3113 -1316 -3111 -1296
rect -3299 -1381 -3297 -1361
rect -3266 -1381 -3264 -1361
rect -3235 -1371 -3233 -1351
rect -122 -1472 -120 -1452
rect -90 -1472 -88 -1452
rect 585 -1470 587 -1430
rect -219 -1496 -217 -1476
rect -167 -1496 -165 -1476
rect -323 -1543 -321 -1523
rect -271 -1543 -269 -1523
rect -219 -1543 -217 -1523
rect -167 -1543 -165 -1523
rect 585 -1535 587 -1495
rect 628 -1504 630 -1484
rect 117 -1640 137 -1638
rect 220 -1652 222 -1632
rect 220 -1685 222 -1665
rect 256 -1687 258 -1667
rect 117 -1691 137 -1689
rect 586 -1753 588 -1713
rect -137 -1809 -135 -1789
rect -105 -1809 -103 -1789
rect 822 -1700 824 -1660
rect 1070 -1657 1072 -1637
rect 1103 -1657 1105 -1637
rect 1134 -1647 1136 -1627
rect 822 -1765 824 -1725
rect 865 -1734 867 -1714
rect -234 -1833 -232 -1813
rect -182 -1833 -180 -1813
rect -338 -1880 -336 -1860
rect -286 -1880 -284 -1860
rect -234 -1880 -232 -1860
rect -182 -1880 -180 -1860
rect 192 -1867 194 -1827
rect 586 -1818 588 -1778
rect 629 -1787 631 -1767
rect 1661 -1681 1681 -1679
rect 1764 -1693 1766 -1673
rect 1764 -1726 1766 -1706
rect 2213 -1678 2215 -1658
rect 2245 -1678 2247 -1658
rect 2116 -1702 2118 -1682
rect 2168 -1702 2170 -1682
rect 1800 -1728 1802 -1708
rect 1661 -1732 1681 -1730
rect 2012 -1749 2014 -1729
rect 2064 -1749 2066 -1729
rect 2116 -1749 2118 -1729
rect 2168 -1749 2170 -1729
rect 1367 -1810 1369 -1790
rect 1400 -1810 1402 -1790
rect 1431 -1800 1433 -1780
rect 192 -1932 194 -1892
rect 235 -1901 237 -1881
rect 831 -1911 833 -1871
rect 582 -2024 584 -1984
rect 831 -1976 833 -1936
rect 874 -1945 876 -1925
rect 1081 -1957 1083 -1937
rect 1114 -1957 1116 -1937
rect 1145 -1947 1147 -1927
rect 582 -2089 584 -2049
rect 625 -2058 627 -2038
rect 570 -2273 572 -2233
rect 570 -2338 572 -2298
rect 613 -2307 615 -2287
rect -137 -2416 -135 -2396
rect -105 -2416 -103 -2396
rect -234 -2440 -232 -2420
rect -182 -2440 -180 -2420
rect -338 -2487 -336 -2467
rect -286 -2487 -284 -2467
rect -234 -2487 -232 -2467
rect -182 -2487 -180 -2467
rect 114 -2515 134 -2513
rect 217 -2527 219 -2507
rect 217 -2560 219 -2540
rect 253 -2562 255 -2542
rect 114 -2566 134 -2564
rect 663 -2620 665 -2580
rect -137 -2686 -135 -2666
rect -105 -2686 -103 -2666
rect -234 -2710 -232 -2690
rect -182 -2710 -180 -2690
rect -338 -2757 -336 -2737
rect -286 -2757 -284 -2737
rect -234 -2757 -232 -2737
rect -182 -2757 -180 -2737
rect 189 -2742 191 -2702
rect 663 -2685 665 -2645
rect 706 -2654 708 -2634
rect 998 -2672 1000 -2632
rect 998 -2737 1000 -2697
rect 1041 -2706 1043 -2686
rect 1294 -2724 1296 -2704
rect 1327 -2724 1329 -2704
rect 1358 -2714 1360 -2694
rect 189 -2807 191 -2767
rect 232 -2776 234 -2756
rect 664 -2903 666 -2863
rect 664 -2968 666 -2928
rect 707 -2937 709 -2917
rect 999 -2955 1001 -2915
rect 999 -3020 1001 -2980
rect 1042 -2989 1044 -2969
rect 2287 -2920 2289 -2900
rect 2319 -2920 2321 -2900
rect 2190 -2944 2192 -2924
rect 2242 -2944 2244 -2924
rect 2086 -2991 2088 -2971
rect 2138 -2991 2140 -2971
rect 2190 -2991 2192 -2971
rect 2242 -2991 2244 -2971
rect 1798 -3038 1800 -3018
rect 1831 -3038 1833 -3018
rect 1862 -3028 1864 -3008
rect 1301 -3113 1303 -3093
rect 1334 -3113 1336 -3093
rect 1365 -3103 1367 -3083
rect 660 -3174 662 -3134
rect 660 -3239 662 -3199
rect 703 -3208 705 -3188
rect 1593 -3269 1595 -3249
rect 1626 -3269 1628 -3249
rect 1657 -3259 1659 -3239
rect 1329 -3357 1331 -3317
rect 648 -3423 650 -3383
rect 648 -3488 650 -3448
rect 691 -3457 693 -3437
rect 1329 -3422 1331 -3382
rect 1372 -3391 1374 -3371
rect 989 -3489 991 -3449
rect 989 -3554 991 -3514
rect 1032 -3523 1034 -3503
rect 665 -3690 667 -3650
rect 665 -3755 667 -3715
rect 708 -3724 710 -3704
rect 653 -3939 655 -3899
rect 653 -4004 655 -3964
rect 696 -3973 698 -3953
<< ptransistor >>
rect 812 1643 852 1645
rect 913 1634 915 1674
rect 1004 1618 1006 1658
rect 1069 1621 1071 1701
rect 1178 1649 1180 1689
rect 1205 1649 1207 1689
rect 812 1592 852 1594
rect 1069 1521 1071 1601
rect 1118 1524 1120 1564
rect 1240 1579 1242 1619
rect 2860 1616 2900 1618
rect 2961 1607 2963 1647
rect 3052 1591 3054 1631
rect 3117 1594 3119 1674
rect 3226 1622 3228 1662
rect 3253 1622 3255 1662
rect 2860 1565 2900 1567
rect 3117 1494 3119 1574
rect 3166 1497 3168 1537
rect 3288 1552 3290 1592
rect -1523 359 -1521 399
rect -1471 359 -1469 399
rect -1419 359 -1417 399
rect -1367 359 -1365 399
rect -1322 367 -1320 407
rect -1290 367 -1288 407
rect 3772 356 3774 396
rect 3824 356 3826 396
rect 3876 356 3878 396
rect 3928 356 3930 396
rect 3973 364 3975 404
rect 4005 364 4007 404
rect -1523 297 -1521 337
rect -1471 297 -1469 337
rect 3772 294 3774 334
rect 3824 294 3826 334
rect 1424 53 1426 93
rect 1476 53 1478 93
rect 1528 53 1530 93
rect 1580 53 1582 93
rect 1625 61 1627 101
rect 1657 61 1659 101
rect -397 -42 -395 -2
rect -345 -42 -343 -2
rect -293 -42 -291 -2
rect -241 -42 -239 -2
rect -196 -34 -194 6
rect -164 -34 -162 6
rect 1071 5 1111 7
rect 1172 -4 1174 36
rect 1424 -9 1426 31
rect 1476 -9 1478 31
rect 1071 -46 1111 -44
rect -397 -104 -395 -64
rect -345 -104 -343 -64
rect 821 -140 823 -60
rect 158 -194 198 -192
rect 259 -203 261 -163
rect 451 -185 453 -145
rect 478 -185 480 -145
rect 158 -245 198 -243
rect -401 -297 -399 -257
rect -349 -297 -347 -257
rect -297 -297 -295 -257
rect -245 -297 -243 -257
rect -200 -289 -198 -249
rect -168 -289 -166 -249
rect 513 -255 515 -215
rect 821 -240 823 -160
rect 870 -237 872 -197
rect 1066 -215 1106 -213
rect 1167 -224 1169 -184
rect 1439 -223 1441 -183
rect 1491 -223 1493 -183
rect 1543 -223 1545 -183
rect 1595 -223 1597 -183
rect 1640 -215 1642 -175
rect 1672 -215 1674 -175
rect -401 -359 -399 -319
rect -349 -359 -347 -319
rect 176 -347 178 -307
rect 203 -347 205 -307
rect 1066 -266 1106 -264
rect 1439 -285 1441 -245
rect 1491 -285 1493 -245
rect 238 -417 240 -377
rect 965 -787 967 -707
rect 1216 -789 1218 -709
rect -304 -879 -302 -839
rect -252 -879 -250 -839
rect -200 -879 -198 -839
rect -148 -879 -146 -839
rect -103 -871 -101 -831
rect -71 -871 -69 -831
rect 631 -836 633 -796
rect 658 -836 660 -796
rect -304 -941 -302 -901
rect -252 -941 -250 -901
rect 693 -906 695 -866
rect 965 -887 967 -807
rect 1014 -884 1016 -844
rect 1216 -889 1218 -809
rect 146 -980 186 -978
rect 247 -989 249 -949
rect 1265 -886 1267 -846
rect 1823 -896 1825 -856
rect 1875 -896 1877 -856
rect 1927 -896 1929 -856
rect 1979 -896 1981 -856
rect 2024 -888 2026 -848
rect 2056 -888 2058 -848
rect 1518 -945 1558 -943
rect 1619 -954 1621 -914
rect 1823 -958 1825 -918
rect 1875 -958 1877 -918
rect 1518 -996 1558 -994
rect 146 -1031 186 -1029
rect -323 -1102 -321 -1062
rect -271 -1102 -269 -1062
rect -219 -1102 -217 -1062
rect -167 -1102 -165 -1062
rect -122 -1094 -120 -1054
rect -90 -1094 -88 -1054
rect 554 -1081 556 -1041
rect 581 -1081 583 -1041
rect 772 -1081 774 -1041
rect 799 -1081 801 -1041
rect -3541 -1214 -3501 -1212
rect -3440 -1223 -3438 -1183
rect -3349 -1239 -3347 -1199
rect -3284 -1236 -3282 -1156
rect -323 -1164 -321 -1124
rect -271 -1164 -269 -1124
rect 164 -1133 166 -1093
rect 191 -1133 193 -1093
rect -3175 -1208 -3173 -1168
rect -3148 -1208 -3146 -1168
rect -3541 -1265 -3501 -1263
rect -3284 -1336 -3282 -1256
rect -3235 -1333 -3233 -1293
rect 226 -1203 228 -1163
rect 616 -1151 618 -1111
rect 834 -1151 836 -1111
rect -3113 -1278 -3111 -1238
rect -323 -1440 -321 -1400
rect -271 -1440 -269 -1400
rect -219 -1440 -217 -1400
rect -167 -1440 -165 -1400
rect -122 -1432 -120 -1392
rect -90 -1432 -88 -1392
rect 566 -1396 568 -1356
rect 593 -1396 595 -1356
rect -323 -1502 -321 -1462
rect -271 -1502 -269 -1462
rect 628 -1466 630 -1426
rect 1085 -1512 1087 -1432
rect 155 -1640 195 -1638
rect 256 -1649 258 -1609
rect 803 -1626 805 -1586
rect 830 -1626 832 -1586
rect 1085 -1612 1087 -1532
rect 567 -1679 569 -1639
rect 594 -1679 596 -1639
rect 1134 -1609 1136 -1569
rect 155 -1691 195 -1689
rect -338 -1777 -336 -1737
rect -286 -1777 -284 -1737
rect -234 -1777 -232 -1737
rect -182 -1777 -180 -1737
rect -137 -1769 -135 -1729
rect -105 -1769 -103 -1729
rect -338 -1839 -336 -1799
rect -286 -1839 -284 -1799
rect 173 -1793 175 -1753
rect 200 -1793 202 -1753
rect 629 -1749 631 -1709
rect 865 -1696 867 -1656
rect 1382 -1665 1384 -1585
rect 2012 -1646 2014 -1606
rect 2064 -1646 2066 -1606
rect 2116 -1646 2118 -1606
rect 2168 -1646 2170 -1606
rect 2213 -1638 2215 -1598
rect 2245 -1638 2247 -1598
rect 235 -1863 237 -1823
rect 812 -1837 814 -1797
rect 839 -1837 841 -1797
rect 1096 -1812 1098 -1732
rect 1382 -1765 1384 -1685
rect 1699 -1681 1739 -1679
rect 1800 -1690 1802 -1650
rect 1431 -1762 1433 -1722
rect 2012 -1708 2014 -1668
rect 2064 -1708 2066 -1668
rect 1699 -1732 1739 -1730
rect 563 -1950 565 -1910
rect 590 -1950 592 -1910
rect 874 -1907 876 -1867
rect 1096 -1912 1098 -1832
rect 1145 -1909 1147 -1869
rect 625 -2020 627 -1980
rect 551 -2199 553 -2159
rect 578 -2199 580 -2159
rect 613 -2269 615 -2229
rect -338 -2384 -336 -2344
rect -286 -2384 -284 -2344
rect -234 -2384 -232 -2344
rect -182 -2384 -180 -2344
rect -137 -2376 -135 -2336
rect -105 -2376 -103 -2336
rect -338 -2446 -336 -2406
rect -286 -2446 -284 -2406
rect 152 -2515 192 -2513
rect 253 -2524 255 -2484
rect 644 -2546 646 -2506
rect 671 -2546 673 -2506
rect 152 -2566 192 -2564
rect -338 -2654 -336 -2614
rect -286 -2654 -284 -2614
rect -234 -2654 -232 -2614
rect -182 -2654 -180 -2614
rect -137 -2646 -135 -2606
rect -105 -2646 -103 -2606
rect -338 -2716 -336 -2676
rect -286 -2716 -284 -2676
rect 170 -2668 172 -2628
rect 197 -2668 199 -2628
rect 706 -2616 708 -2576
rect 979 -2598 981 -2558
rect 1006 -2598 1008 -2558
rect 1309 -2579 1311 -2499
rect 1041 -2668 1043 -2628
rect 1309 -2679 1311 -2599
rect 232 -2738 234 -2698
rect 1358 -2676 1360 -2636
rect 645 -2829 647 -2789
rect 672 -2829 674 -2789
rect 707 -2899 709 -2859
rect 980 -2881 982 -2841
rect 1007 -2881 1009 -2841
rect 1042 -2951 1044 -2911
rect 1316 -2968 1318 -2888
rect 1813 -2893 1815 -2813
rect 2086 -2888 2088 -2848
rect 2138 -2888 2140 -2848
rect 2190 -2888 2192 -2848
rect 2242 -2888 2244 -2848
rect 2287 -2880 2289 -2840
rect 2319 -2880 2321 -2840
rect 641 -3100 643 -3060
rect 668 -3100 670 -3060
rect 1316 -3068 1318 -2988
rect 1813 -2993 1815 -2913
rect 2086 -2950 2088 -2910
rect 2138 -2950 2140 -2910
rect 1862 -2990 1864 -2950
rect 1365 -3065 1367 -3025
rect 1608 -3124 1610 -3044
rect 703 -3170 705 -3130
rect 1608 -3224 1610 -3144
rect 1310 -3283 1312 -3243
rect 1337 -3283 1339 -3243
rect 1657 -3221 1659 -3181
rect 629 -3349 631 -3309
rect 656 -3349 658 -3309
rect 1372 -3353 1374 -3313
rect 691 -3419 693 -3379
rect 970 -3415 972 -3375
rect 997 -3415 999 -3375
rect 1032 -3485 1034 -3445
rect 646 -3616 648 -3576
rect 673 -3616 675 -3576
rect 708 -3686 710 -3646
rect 634 -3865 636 -3825
rect 661 -3865 663 -3825
rect 696 -3935 698 -3895
<< ndiffusion >>
rect 774 1645 794 1646
rect 774 1642 794 1643
rect 876 1631 877 1651
rect 879 1631 880 1651
rect 774 1594 794 1595
rect 876 1598 877 1618
rect 879 1598 880 1618
rect 912 1596 913 1616
rect 915 1596 916 1616
rect 774 1591 794 1592
rect 1003 1580 1004 1600
rect 1006 1580 1007 1600
rect 1196 1575 1197 1615
rect 1199 1575 1200 1615
rect 2822 1618 2842 1619
rect 2822 1615 2842 1616
rect 2924 1604 2925 1624
rect 2927 1604 2928 1624
rect 2822 1567 2842 1568
rect 2924 1571 2925 1591
rect 2927 1571 2928 1591
rect 2960 1569 2961 1589
rect 2963 1569 2964 1589
rect 2822 1564 2842 1565
rect 1196 1510 1197 1550
rect 1199 1510 1200 1550
rect 1239 1541 1240 1561
rect 1242 1541 1243 1561
rect 3051 1553 3052 1573
rect 3054 1553 3055 1573
rect 1053 1476 1054 1496
rect 1056 1476 1057 1496
rect 1086 1476 1087 1496
rect 1089 1476 1090 1496
rect 1117 1486 1118 1506
rect 1120 1486 1121 1506
rect 3244 1548 3245 1588
rect 3247 1548 3248 1588
rect 3244 1483 3245 1523
rect 3247 1483 3248 1523
rect 3287 1514 3288 1534
rect 3290 1514 3291 1534
rect 3101 1449 3102 1469
rect 3104 1449 3105 1469
rect 3134 1449 3135 1469
rect 3137 1449 3138 1469
rect 3165 1459 3166 1479
rect 3168 1459 3169 1479
rect -1323 327 -1322 347
rect -1320 327 -1319 347
rect -1291 327 -1290 347
rect -1288 327 -1287 347
rect -1420 303 -1419 323
rect -1417 303 -1416 323
rect -1368 303 -1367 323
rect -1365 303 -1364 323
rect 3972 324 3973 344
rect 3975 324 3976 344
rect 4004 324 4005 344
rect 4007 324 4008 344
rect 3875 300 3876 320
rect 3878 300 3879 320
rect 3927 300 3928 320
rect 3930 300 3931 320
rect -1524 256 -1523 276
rect -1521 256 -1520 276
rect -1472 256 -1471 276
rect -1469 256 -1468 276
rect -1420 256 -1419 276
rect -1417 256 -1416 276
rect -1368 256 -1367 276
rect -1365 256 -1364 276
rect 3771 253 3772 273
rect 3774 253 3775 273
rect 3823 253 3824 273
rect 3826 253 3827 273
rect 3875 253 3876 273
rect 3878 253 3879 273
rect 3927 253 3928 273
rect 3930 253 3931 273
rect 1033 7 1053 8
rect 1033 4 1053 5
rect 1135 -7 1136 13
rect 1138 -7 1139 13
rect 1033 -44 1053 -43
rect 1135 -40 1136 -20
rect 1138 -40 1139 -20
rect 1624 21 1625 41
rect 1627 21 1628 41
rect 1656 21 1657 41
rect 1659 21 1660 41
rect 1527 -3 1528 17
rect 1530 -3 1531 17
rect 1579 -3 1580 17
rect 1582 -3 1583 17
rect 1171 -42 1172 -22
rect 1174 -42 1175 -22
rect 1033 -47 1053 -46
rect -197 -74 -196 -54
rect -194 -74 -193 -54
rect -165 -74 -164 -54
rect -162 -74 -161 -54
rect 1423 -50 1424 -30
rect 1426 -50 1427 -30
rect 1475 -50 1476 -30
rect 1478 -50 1479 -30
rect 1527 -50 1528 -30
rect 1530 -50 1531 -30
rect 1579 -50 1580 -30
rect 1582 -50 1583 -30
rect -294 -98 -293 -78
rect -291 -98 -290 -78
rect -242 -98 -241 -78
rect -239 -98 -238 -78
rect -398 -145 -397 -125
rect -395 -145 -394 -125
rect -346 -145 -345 -125
rect -343 -145 -342 -125
rect -294 -145 -293 -125
rect -291 -145 -290 -125
rect -242 -145 -241 -125
rect -239 -145 -238 -125
rect 120 -192 140 -191
rect 120 -195 140 -194
rect 222 -206 223 -186
rect 225 -206 226 -186
rect 120 -243 140 -242
rect 222 -239 223 -219
rect 225 -239 226 -219
rect 258 -241 259 -221
rect 261 -241 262 -221
rect 120 -246 140 -245
rect 469 -259 470 -219
rect 472 -259 473 -219
rect 1028 -213 1048 -212
rect 1028 -216 1048 -215
rect 1130 -227 1131 -207
rect 1133 -227 1134 -207
rect -201 -329 -200 -309
rect -198 -329 -197 -309
rect -169 -329 -168 -309
rect -166 -329 -165 -309
rect -298 -353 -297 -333
rect -295 -353 -294 -333
rect -246 -353 -245 -333
rect -243 -353 -242 -333
rect 469 -324 470 -284
rect 472 -324 473 -284
rect 512 -293 513 -273
rect 515 -293 516 -273
rect 805 -285 806 -265
rect 808 -285 809 -265
rect 838 -285 839 -265
rect 841 -285 842 -265
rect 869 -275 870 -255
rect 872 -275 873 -255
rect 1028 -264 1048 -263
rect 1130 -260 1131 -240
rect 1133 -260 1134 -240
rect 1166 -262 1167 -242
rect 1169 -262 1170 -242
rect 1028 -267 1048 -266
rect 1639 -255 1640 -235
rect 1642 -255 1643 -235
rect 1671 -255 1672 -235
rect 1674 -255 1675 -235
rect 1542 -279 1543 -259
rect 1545 -279 1546 -259
rect 1594 -279 1595 -259
rect 1597 -279 1598 -259
rect 1438 -326 1439 -306
rect 1441 -326 1442 -306
rect 1490 -326 1491 -306
rect 1493 -326 1494 -306
rect 1542 -326 1543 -306
rect 1545 -326 1546 -306
rect 1594 -326 1595 -306
rect 1597 -326 1598 -306
rect -402 -400 -401 -380
rect -399 -400 -398 -380
rect -350 -400 -349 -380
rect -347 -400 -346 -380
rect -298 -400 -297 -380
rect -295 -400 -294 -380
rect -246 -400 -245 -380
rect -243 -400 -242 -380
rect 194 -421 195 -381
rect 197 -421 198 -381
rect 194 -486 195 -446
rect 197 -486 198 -446
rect 237 -455 238 -435
rect 240 -455 241 -435
rect -104 -911 -103 -891
rect -101 -911 -100 -891
rect -72 -911 -71 -891
rect -69 -911 -68 -891
rect 649 -910 650 -870
rect 652 -910 653 -870
rect -201 -935 -200 -915
rect -198 -935 -197 -915
rect -149 -935 -148 -915
rect -146 -935 -145 -915
rect -305 -982 -304 -962
rect -302 -982 -301 -962
rect -253 -982 -252 -962
rect -250 -982 -249 -962
rect -201 -982 -200 -962
rect -198 -982 -197 -962
rect -149 -982 -148 -962
rect -146 -982 -145 -962
rect 108 -978 128 -977
rect 108 -981 128 -980
rect 210 -992 211 -972
rect 213 -992 214 -972
rect 649 -975 650 -935
rect 652 -975 653 -935
rect 692 -944 693 -924
rect 695 -944 696 -924
rect 949 -932 950 -912
rect 952 -932 953 -912
rect 982 -932 983 -912
rect 985 -932 986 -912
rect 1013 -922 1014 -902
rect 1016 -922 1017 -902
rect 1200 -934 1201 -914
rect 1203 -934 1204 -914
rect 1233 -934 1234 -914
rect 1236 -934 1237 -914
rect 1264 -924 1265 -904
rect 1267 -924 1268 -904
rect 1480 -943 1500 -942
rect 1480 -946 1500 -945
rect 1582 -957 1583 -937
rect 1585 -957 1586 -937
rect 108 -1029 128 -1028
rect 210 -1025 211 -1005
rect 213 -1025 214 -1005
rect 1480 -994 1500 -993
rect 1582 -990 1583 -970
rect 1585 -990 1586 -970
rect 2023 -928 2024 -908
rect 2026 -928 2027 -908
rect 2055 -928 2056 -908
rect 2058 -928 2059 -908
rect 1926 -952 1927 -932
rect 1929 -952 1930 -932
rect 1978 -952 1979 -932
rect 1981 -952 1982 -932
rect 1618 -992 1619 -972
rect 1621 -992 1622 -972
rect 1480 -997 1500 -996
rect 1822 -999 1823 -979
rect 1825 -999 1826 -979
rect 1874 -999 1875 -979
rect 1877 -999 1878 -979
rect 1926 -999 1927 -979
rect 1929 -999 1930 -979
rect 1978 -999 1979 -979
rect 1981 -999 1982 -979
rect 246 -1027 247 -1007
rect 249 -1027 250 -1007
rect 108 -1032 128 -1031
rect -3579 -1212 -3559 -1211
rect -3579 -1215 -3559 -1214
rect -3477 -1226 -3476 -1206
rect -3474 -1226 -3473 -1206
rect -3579 -1263 -3559 -1262
rect -3477 -1259 -3476 -1239
rect -3474 -1259 -3473 -1239
rect -123 -1134 -122 -1114
rect -120 -1134 -119 -1114
rect -91 -1134 -90 -1114
rect -88 -1134 -87 -1114
rect -220 -1158 -219 -1138
rect -217 -1158 -216 -1138
rect -168 -1158 -167 -1138
rect -165 -1158 -164 -1138
rect -324 -1205 -323 -1185
rect -321 -1205 -320 -1185
rect -272 -1205 -271 -1185
rect -269 -1205 -268 -1185
rect -220 -1205 -219 -1185
rect -217 -1205 -216 -1185
rect -168 -1205 -167 -1185
rect -165 -1205 -164 -1185
rect -3441 -1261 -3440 -1241
rect -3438 -1261 -3437 -1241
rect 182 -1207 183 -1167
rect 185 -1207 186 -1167
rect -3579 -1266 -3559 -1265
rect -3350 -1277 -3349 -1257
rect -3347 -1277 -3346 -1257
rect -3157 -1282 -3156 -1242
rect -3154 -1282 -3153 -1242
rect 572 -1155 573 -1115
rect 575 -1155 576 -1115
rect 790 -1155 791 -1115
rect 793 -1155 794 -1115
rect 572 -1220 573 -1180
rect 575 -1220 576 -1180
rect 615 -1189 616 -1169
rect 618 -1189 619 -1169
rect 790 -1220 791 -1180
rect 793 -1220 794 -1180
rect 833 -1189 834 -1169
rect 836 -1189 837 -1169
rect 182 -1272 183 -1232
rect 185 -1272 186 -1232
rect 225 -1241 226 -1221
rect 228 -1241 229 -1221
rect -3157 -1347 -3156 -1307
rect -3154 -1347 -3153 -1307
rect -3114 -1316 -3113 -1296
rect -3111 -1316 -3110 -1296
rect -3300 -1381 -3299 -1361
rect -3297 -1381 -3296 -1361
rect -3267 -1381 -3266 -1361
rect -3264 -1381 -3263 -1361
rect -3236 -1371 -3235 -1351
rect -3233 -1371 -3232 -1351
rect -123 -1472 -122 -1452
rect -120 -1472 -119 -1452
rect -91 -1472 -90 -1452
rect -88 -1472 -87 -1452
rect 584 -1470 585 -1430
rect 587 -1470 588 -1430
rect -220 -1496 -219 -1476
rect -217 -1496 -216 -1476
rect -168 -1496 -167 -1476
rect -165 -1496 -164 -1476
rect -324 -1543 -323 -1523
rect -321 -1543 -320 -1523
rect -272 -1543 -271 -1523
rect -269 -1543 -268 -1523
rect -220 -1543 -219 -1523
rect -217 -1543 -216 -1523
rect -168 -1543 -167 -1523
rect -165 -1543 -164 -1523
rect 584 -1535 585 -1495
rect 587 -1535 588 -1495
rect 627 -1504 628 -1484
rect 630 -1504 631 -1484
rect 117 -1638 137 -1637
rect 117 -1641 137 -1640
rect 219 -1652 220 -1632
rect 222 -1652 223 -1632
rect 117 -1689 137 -1688
rect 219 -1685 220 -1665
rect 222 -1685 223 -1665
rect 255 -1687 256 -1667
rect 258 -1687 259 -1667
rect 117 -1692 137 -1691
rect 585 -1753 586 -1713
rect 588 -1753 589 -1713
rect -138 -1809 -137 -1789
rect -135 -1809 -134 -1789
rect -106 -1809 -105 -1789
rect -103 -1809 -102 -1789
rect 821 -1700 822 -1660
rect 824 -1700 825 -1660
rect 1069 -1657 1070 -1637
rect 1072 -1657 1073 -1637
rect 1102 -1657 1103 -1637
rect 1105 -1657 1106 -1637
rect 1133 -1647 1134 -1627
rect 1136 -1647 1137 -1627
rect 821 -1765 822 -1725
rect 824 -1765 825 -1725
rect 864 -1734 865 -1714
rect 867 -1734 868 -1714
rect -235 -1833 -234 -1813
rect -232 -1833 -231 -1813
rect -183 -1833 -182 -1813
rect -180 -1833 -179 -1813
rect -339 -1880 -338 -1860
rect -336 -1880 -335 -1860
rect -287 -1880 -286 -1860
rect -284 -1880 -283 -1860
rect -235 -1880 -234 -1860
rect -232 -1880 -231 -1860
rect -183 -1880 -182 -1860
rect -180 -1880 -179 -1860
rect 191 -1867 192 -1827
rect 194 -1867 195 -1827
rect 585 -1818 586 -1778
rect 588 -1818 589 -1778
rect 628 -1787 629 -1767
rect 631 -1787 632 -1767
rect 1661 -1679 1681 -1678
rect 1661 -1682 1681 -1681
rect 1763 -1693 1764 -1673
rect 1766 -1693 1767 -1673
rect 1661 -1730 1681 -1729
rect 1763 -1726 1764 -1706
rect 1766 -1726 1767 -1706
rect 2212 -1678 2213 -1658
rect 2215 -1678 2216 -1658
rect 2244 -1678 2245 -1658
rect 2247 -1678 2248 -1658
rect 2115 -1702 2116 -1682
rect 2118 -1702 2119 -1682
rect 2167 -1702 2168 -1682
rect 2170 -1702 2171 -1682
rect 1799 -1728 1800 -1708
rect 1802 -1728 1803 -1708
rect 1661 -1733 1681 -1732
rect 2011 -1749 2012 -1729
rect 2014 -1749 2015 -1729
rect 2063 -1749 2064 -1729
rect 2066 -1749 2067 -1729
rect 2115 -1749 2116 -1729
rect 2118 -1749 2119 -1729
rect 2167 -1749 2168 -1729
rect 2170 -1749 2171 -1729
rect 1366 -1810 1367 -1790
rect 1369 -1810 1370 -1790
rect 1399 -1810 1400 -1790
rect 1402 -1810 1403 -1790
rect 1430 -1800 1431 -1780
rect 1433 -1800 1434 -1780
rect 191 -1932 192 -1892
rect 194 -1932 195 -1892
rect 234 -1901 235 -1881
rect 237 -1901 238 -1881
rect 830 -1911 831 -1871
rect 833 -1911 834 -1871
rect 581 -2024 582 -1984
rect 584 -2024 585 -1984
rect 830 -1976 831 -1936
rect 833 -1976 834 -1936
rect 873 -1945 874 -1925
rect 876 -1945 877 -1925
rect 1080 -1957 1081 -1937
rect 1083 -1957 1084 -1937
rect 1113 -1957 1114 -1937
rect 1116 -1957 1117 -1937
rect 1144 -1947 1145 -1927
rect 1147 -1947 1148 -1927
rect 581 -2089 582 -2049
rect 584 -2089 585 -2049
rect 624 -2058 625 -2038
rect 627 -2058 628 -2038
rect 569 -2273 570 -2233
rect 572 -2273 573 -2233
rect 569 -2338 570 -2298
rect 572 -2338 573 -2298
rect 612 -2307 613 -2287
rect 615 -2307 616 -2287
rect -138 -2416 -137 -2396
rect -135 -2416 -134 -2396
rect -106 -2416 -105 -2396
rect -103 -2416 -102 -2396
rect -235 -2440 -234 -2420
rect -232 -2440 -231 -2420
rect -183 -2440 -182 -2420
rect -180 -2440 -179 -2420
rect -339 -2487 -338 -2467
rect -336 -2487 -335 -2467
rect -287 -2487 -286 -2467
rect -284 -2487 -283 -2467
rect -235 -2487 -234 -2467
rect -232 -2487 -231 -2467
rect -183 -2487 -182 -2467
rect -180 -2487 -179 -2467
rect 114 -2513 134 -2512
rect 114 -2516 134 -2515
rect 216 -2527 217 -2507
rect 219 -2527 220 -2507
rect 114 -2564 134 -2563
rect 216 -2560 217 -2540
rect 219 -2560 220 -2540
rect 252 -2562 253 -2542
rect 255 -2562 256 -2542
rect 114 -2567 134 -2566
rect 662 -2620 663 -2580
rect 665 -2620 666 -2580
rect -138 -2686 -137 -2666
rect -135 -2686 -134 -2666
rect -106 -2686 -105 -2666
rect -103 -2686 -102 -2666
rect -235 -2710 -234 -2690
rect -232 -2710 -231 -2690
rect -183 -2710 -182 -2690
rect -180 -2710 -179 -2690
rect -339 -2757 -338 -2737
rect -336 -2757 -335 -2737
rect -287 -2757 -286 -2737
rect -284 -2757 -283 -2737
rect -235 -2757 -234 -2737
rect -232 -2757 -231 -2737
rect -183 -2757 -182 -2737
rect -180 -2757 -179 -2737
rect 188 -2742 189 -2702
rect 191 -2742 192 -2702
rect 662 -2685 663 -2645
rect 665 -2685 666 -2645
rect 705 -2654 706 -2634
rect 708 -2654 709 -2634
rect 997 -2672 998 -2632
rect 1000 -2672 1001 -2632
rect 997 -2737 998 -2697
rect 1000 -2737 1001 -2697
rect 1040 -2706 1041 -2686
rect 1043 -2706 1044 -2686
rect 1293 -2724 1294 -2704
rect 1296 -2724 1297 -2704
rect 1326 -2724 1327 -2704
rect 1329 -2724 1330 -2704
rect 1357 -2714 1358 -2694
rect 1360 -2714 1361 -2694
rect 188 -2807 189 -2767
rect 191 -2807 192 -2767
rect 231 -2776 232 -2756
rect 234 -2776 235 -2756
rect 663 -2903 664 -2863
rect 666 -2903 667 -2863
rect 663 -2968 664 -2928
rect 666 -2968 667 -2928
rect 706 -2937 707 -2917
rect 709 -2937 710 -2917
rect 998 -2955 999 -2915
rect 1001 -2955 1002 -2915
rect 998 -3020 999 -2980
rect 1001 -3020 1002 -2980
rect 1041 -2989 1042 -2969
rect 1044 -2989 1045 -2969
rect 2286 -2920 2287 -2900
rect 2289 -2920 2290 -2900
rect 2318 -2920 2319 -2900
rect 2321 -2920 2322 -2900
rect 2189 -2944 2190 -2924
rect 2192 -2944 2193 -2924
rect 2241 -2944 2242 -2924
rect 2244 -2944 2245 -2924
rect 2085 -2991 2086 -2971
rect 2088 -2991 2089 -2971
rect 2137 -2991 2138 -2971
rect 2140 -2991 2141 -2971
rect 2189 -2991 2190 -2971
rect 2192 -2991 2193 -2971
rect 2241 -2991 2242 -2971
rect 2244 -2991 2245 -2971
rect 1797 -3038 1798 -3018
rect 1800 -3038 1801 -3018
rect 1830 -3038 1831 -3018
rect 1833 -3038 1834 -3018
rect 1861 -3028 1862 -3008
rect 1864 -3028 1865 -3008
rect 1300 -3113 1301 -3093
rect 1303 -3113 1304 -3093
rect 1333 -3113 1334 -3093
rect 1336 -3113 1337 -3093
rect 1364 -3103 1365 -3083
rect 1367 -3103 1368 -3083
rect 659 -3174 660 -3134
rect 662 -3174 663 -3134
rect 659 -3239 660 -3199
rect 662 -3239 663 -3199
rect 702 -3208 703 -3188
rect 705 -3208 706 -3188
rect 1592 -3269 1593 -3249
rect 1595 -3269 1596 -3249
rect 1625 -3269 1626 -3249
rect 1628 -3269 1629 -3249
rect 1656 -3259 1657 -3239
rect 1659 -3259 1660 -3239
rect 1328 -3357 1329 -3317
rect 1331 -3357 1332 -3317
rect 647 -3423 648 -3383
rect 650 -3423 651 -3383
rect 647 -3488 648 -3448
rect 650 -3488 651 -3448
rect 690 -3457 691 -3437
rect 693 -3457 694 -3437
rect 1328 -3422 1329 -3382
rect 1331 -3422 1332 -3382
rect 1371 -3391 1372 -3371
rect 1374 -3391 1375 -3371
rect 988 -3489 989 -3449
rect 991 -3489 992 -3449
rect 988 -3554 989 -3514
rect 991 -3554 992 -3514
rect 1031 -3523 1032 -3503
rect 1034 -3523 1035 -3503
rect 664 -3690 665 -3650
rect 667 -3690 668 -3650
rect 664 -3755 665 -3715
rect 667 -3755 668 -3715
rect 707 -3724 708 -3704
rect 710 -3724 711 -3704
rect 652 -3939 653 -3899
rect 655 -3939 656 -3899
rect 652 -4004 653 -3964
rect 655 -4004 656 -3964
rect 695 -3973 696 -3953
rect 698 -3973 699 -3953
<< pdiffusion >>
rect 812 1645 852 1646
rect 812 1642 852 1643
rect 912 1634 913 1674
rect 915 1634 916 1674
rect 1003 1618 1004 1658
rect 1006 1618 1007 1658
rect 1068 1621 1069 1701
rect 1071 1621 1072 1701
rect 1177 1649 1178 1689
rect 1180 1649 1181 1689
rect 1204 1649 1205 1689
rect 1207 1649 1208 1689
rect 812 1594 852 1595
rect 812 1591 852 1592
rect 1068 1521 1069 1601
rect 1071 1521 1072 1601
rect 1117 1524 1118 1564
rect 1120 1524 1121 1564
rect 1239 1579 1240 1619
rect 1242 1579 1243 1619
rect 2860 1618 2900 1619
rect 2860 1615 2900 1616
rect 2960 1607 2961 1647
rect 2963 1607 2964 1647
rect 3051 1591 3052 1631
rect 3054 1591 3055 1631
rect 3116 1594 3117 1674
rect 3119 1594 3120 1674
rect 3225 1622 3226 1662
rect 3228 1622 3229 1662
rect 3252 1622 3253 1662
rect 3255 1622 3256 1662
rect 2860 1567 2900 1568
rect 2860 1564 2900 1565
rect 3116 1494 3117 1574
rect 3119 1494 3120 1574
rect 3165 1497 3166 1537
rect 3168 1497 3169 1537
rect 3287 1552 3288 1592
rect 3290 1552 3291 1592
rect -1524 359 -1523 399
rect -1521 359 -1520 399
rect -1472 359 -1471 399
rect -1469 359 -1468 399
rect -1420 359 -1419 399
rect -1417 359 -1416 399
rect -1368 359 -1367 399
rect -1365 359 -1364 399
rect -1323 367 -1322 407
rect -1320 367 -1319 407
rect -1291 367 -1290 407
rect -1288 367 -1287 407
rect 3771 356 3772 396
rect 3774 356 3775 396
rect 3823 356 3824 396
rect 3826 356 3827 396
rect 3875 356 3876 396
rect 3878 356 3879 396
rect 3927 356 3928 396
rect 3930 356 3931 396
rect 3972 364 3973 404
rect 3975 364 3976 404
rect 4004 364 4005 404
rect 4007 364 4008 404
rect -1524 297 -1523 337
rect -1521 297 -1520 337
rect -1472 297 -1471 337
rect -1469 297 -1468 337
rect 3771 294 3772 334
rect 3774 294 3775 334
rect 3823 294 3824 334
rect 3826 294 3827 334
rect 1423 53 1424 93
rect 1426 53 1427 93
rect 1475 53 1476 93
rect 1478 53 1479 93
rect 1527 53 1528 93
rect 1530 53 1531 93
rect 1579 53 1580 93
rect 1582 53 1583 93
rect 1624 61 1625 101
rect 1627 61 1628 101
rect 1656 61 1657 101
rect 1659 61 1660 101
rect 1071 7 1111 8
rect -398 -42 -397 -2
rect -395 -42 -394 -2
rect -346 -42 -345 -2
rect -343 -42 -342 -2
rect -294 -42 -293 -2
rect -291 -42 -290 -2
rect -242 -42 -241 -2
rect -239 -42 -238 -2
rect -197 -34 -196 6
rect -194 -34 -193 6
rect -165 -34 -164 6
rect -162 -34 -161 6
rect 1071 4 1111 5
rect 1171 -4 1172 36
rect 1174 -4 1175 36
rect 1423 -9 1424 31
rect 1426 -9 1427 31
rect 1475 -9 1476 31
rect 1478 -9 1479 31
rect 1071 -44 1111 -43
rect 1071 -47 1111 -46
rect -398 -104 -397 -64
rect -395 -104 -394 -64
rect -346 -104 -345 -64
rect -343 -104 -342 -64
rect 820 -140 821 -60
rect 823 -140 824 -60
rect 158 -192 198 -191
rect 158 -195 198 -194
rect 258 -203 259 -163
rect 261 -203 262 -163
rect 450 -185 451 -145
rect 453 -185 454 -145
rect 477 -185 478 -145
rect 480 -185 481 -145
rect 158 -243 198 -242
rect -402 -297 -401 -257
rect -399 -297 -398 -257
rect -350 -297 -349 -257
rect -347 -297 -346 -257
rect -298 -297 -297 -257
rect -295 -297 -294 -257
rect -246 -297 -245 -257
rect -243 -297 -242 -257
rect -201 -289 -200 -249
rect -198 -289 -197 -249
rect -169 -289 -168 -249
rect -166 -289 -165 -249
rect 158 -246 198 -245
rect 512 -255 513 -215
rect 515 -255 516 -215
rect 820 -240 821 -160
rect 823 -240 824 -160
rect 869 -237 870 -197
rect 872 -237 873 -197
rect 1066 -213 1106 -212
rect 1066 -216 1106 -215
rect 1166 -224 1167 -184
rect 1169 -224 1170 -184
rect 1438 -223 1439 -183
rect 1441 -223 1442 -183
rect 1490 -223 1491 -183
rect 1493 -223 1494 -183
rect 1542 -223 1543 -183
rect 1545 -223 1546 -183
rect 1594 -223 1595 -183
rect 1597 -223 1598 -183
rect 1639 -215 1640 -175
rect 1642 -215 1643 -175
rect 1671 -215 1672 -175
rect 1674 -215 1675 -175
rect -402 -359 -401 -319
rect -399 -359 -398 -319
rect -350 -359 -349 -319
rect -347 -359 -346 -319
rect 175 -347 176 -307
rect 178 -347 179 -307
rect 202 -347 203 -307
rect 205 -347 206 -307
rect 1066 -264 1106 -263
rect 1066 -267 1106 -266
rect 1438 -285 1439 -245
rect 1441 -285 1442 -245
rect 1490 -285 1491 -245
rect 1493 -285 1494 -245
rect 237 -417 238 -377
rect 240 -417 241 -377
rect 964 -787 965 -707
rect 967 -787 968 -707
rect 1215 -789 1216 -709
rect 1218 -789 1219 -709
rect -305 -879 -304 -839
rect -302 -879 -301 -839
rect -253 -879 -252 -839
rect -250 -879 -249 -839
rect -201 -879 -200 -839
rect -198 -879 -197 -839
rect -149 -879 -148 -839
rect -146 -879 -145 -839
rect -104 -871 -103 -831
rect -101 -871 -100 -831
rect -72 -871 -71 -831
rect -69 -871 -68 -831
rect 630 -836 631 -796
rect 633 -836 634 -796
rect 657 -836 658 -796
rect 660 -836 661 -796
rect -305 -941 -304 -901
rect -302 -941 -301 -901
rect -253 -941 -252 -901
rect -250 -941 -249 -901
rect 692 -906 693 -866
rect 695 -906 696 -866
rect 964 -887 965 -807
rect 967 -887 968 -807
rect 1013 -884 1014 -844
rect 1016 -884 1017 -844
rect 1215 -889 1216 -809
rect 1218 -889 1219 -809
rect 146 -978 186 -977
rect 146 -981 186 -980
rect 246 -989 247 -949
rect 249 -989 250 -949
rect 1264 -886 1265 -846
rect 1267 -886 1268 -846
rect 1822 -896 1823 -856
rect 1825 -896 1826 -856
rect 1874 -896 1875 -856
rect 1877 -896 1878 -856
rect 1926 -896 1927 -856
rect 1929 -896 1930 -856
rect 1978 -896 1979 -856
rect 1981 -896 1982 -856
rect 2023 -888 2024 -848
rect 2026 -888 2027 -848
rect 2055 -888 2056 -848
rect 2058 -888 2059 -848
rect 1518 -943 1558 -942
rect 1518 -946 1558 -945
rect 1618 -954 1619 -914
rect 1621 -954 1622 -914
rect 1822 -958 1823 -918
rect 1825 -958 1826 -918
rect 1874 -958 1875 -918
rect 1877 -958 1878 -918
rect 1518 -994 1558 -993
rect 1518 -997 1558 -996
rect 146 -1029 186 -1028
rect 146 -1032 186 -1031
rect -324 -1102 -323 -1062
rect -321 -1102 -320 -1062
rect -272 -1102 -271 -1062
rect -269 -1102 -268 -1062
rect -220 -1102 -219 -1062
rect -217 -1102 -216 -1062
rect -168 -1102 -167 -1062
rect -165 -1102 -164 -1062
rect -123 -1094 -122 -1054
rect -120 -1094 -119 -1054
rect -91 -1094 -90 -1054
rect -88 -1094 -87 -1054
rect 553 -1081 554 -1041
rect 556 -1081 557 -1041
rect 580 -1081 581 -1041
rect 583 -1081 584 -1041
rect 771 -1081 772 -1041
rect 774 -1081 775 -1041
rect 798 -1081 799 -1041
rect 801 -1081 802 -1041
rect -3541 -1212 -3501 -1211
rect -3541 -1215 -3501 -1214
rect -3441 -1223 -3440 -1183
rect -3438 -1223 -3437 -1183
rect -3350 -1239 -3349 -1199
rect -3347 -1239 -3346 -1199
rect -3285 -1236 -3284 -1156
rect -3282 -1236 -3281 -1156
rect -324 -1164 -323 -1124
rect -321 -1164 -320 -1124
rect -272 -1164 -271 -1124
rect -269 -1164 -268 -1124
rect 163 -1133 164 -1093
rect 166 -1133 167 -1093
rect 190 -1133 191 -1093
rect 193 -1133 194 -1093
rect -3176 -1208 -3175 -1168
rect -3173 -1208 -3172 -1168
rect -3149 -1208 -3148 -1168
rect -3146 -1208 -3145 -1168
rect -3541 -1263 -3501 -1262
rect -3541 -1266 -3501 -1265
rect -3285 -1336 -3284 -1256
rect -3282 -1336 -3281 -1256
rect -3236 -1333 -3235 -1293
rect -3233 -1333 -3232 -1293
rect 225 -1203 226 -1163
rect 228 -1203 229 -1163
rect 615 -1151 616 -1111
rect 618 -1151 619 -1111
rect 833 -1151 834 -1111
rect 836 -1151 837 -1111
rect -3114 -1278 -3113 -1238
rect -3111 -1278 -3110 -1238
rect -324 -1440 -323 -1400
rect -321 -1440 -320 -1400
rect -272 -1440 -271 -1400
rect -269 -1440 -268 -1400
rect -220 -1440 -219 -1400
rect -217 -1440 -216 -1400
rect -168 -1440 -167 -1400
rect -165 -1440 -164 -1400
rect -123 -1432 -122 -1392
rect -120 -1432 -119 -1392
rect -91 -1432 -90 -1392
rect -88 -1432 -87 -1392
rect 565 -1396 566 -1356
rect 568 -1396 569 -1356
rect 592 -1396 593 -1356
rect 595 -1396 596 -1356
rect -324 -1502 -323 -1462
rect -321 -1502 -320 -1462
rect -272 -1502 -271 -1462
rect -269 -1502 -268 -1462
rect 627 -1466 628 -1426
rect 630 -1466 631 -1426
rect 1084 -1512 1085 -1432
rect 1087 -1512 1088 -1432
rect 155 -1638 195 -1637
rect 155 -1641 195 -1640
rect 255 -1649 256 -1609
rect 258 -1649 259 -1609
rect 802 -1626 803 -1586
rect 805 -1626 806 -1586
rect 829 -1626 830 -1586
rect 832 -1626 833 -1586
rect 1084 -1612 1085 -1532
rect 1087 -1612 1088 -1532
rect 566 -1679 567 -1639
rect 569 -1679 570 -1639
rect 593 -1679 594 -1639
rect 596 -1679 597 -1639
rect 1133 -1609 1134 -1569
rect 1136 -1609 1137 -1569
rect 155 -1689 195 -1688
rect 155 -1692 195 -1691
rect -339 -1777 -338 -1737
rect -336 -1777 -335 -1737
rect -287 -1777 -286 -1737
rect -284 -1777 -283 -1737
rect -235 -1777 -234 -1737
rect -232 -1777 -231 -1737
rect -183 -1777 -182 -1737
rect -180 -1777 -179 -1737
rect -138 -1769 -137 -1729
rect -135 -1769 -134 -1729
rect -106 -1769 -105 -1729
rect -103 -1769 -102 -1729
rect -339 -1839 -338 -1799
rect -336 -1839 -335 -1799
rect -287 -1839 -286 -1799
rect -284 -1839 -283 -1799
rect 172 -1793 173 -1753
rect 175 -1793 176 -1753
rect 199 -1793 200 -1753
rect 202 -1793 203 -1753
rect 628 -1749 629 -1709
rect 631 -1749 632 -1709
rect 864 -1696 865 -1656
rect 867 -1696 868 -1656
rect 1381 -1665 1382 -1585
rect 1384 -1665 1385 -1585
rect 2011 -1646 2012 -1606
rect 2014 -1646 2015 -1606
rect 2063 -1646 2064 -1606
rect 2066 -1646 2067 -1606
rect 2115 -1646 2116 -1606
rect 2118 -1646 2119 -1606
rect 2167 -1646 2168 -1606
rect 2170 -1646 2171 -1606
rect 2212 -1638 2213 -1598
rect 2215 -1638 2216 -1598
rect 2244 -1638 2245 -1598
rect 2247 -1638 2248 -1598
rect 234 -1863 235 -1823
rect 237 -1863 238 -1823
rect 811 -1837 812 -1797
rect 814 -1837 815 -1797
rect 838 -1837 839 -1797
rect 841 -1837 842 -1797
rect 1095 -1812 1096 -1732
rect 1098 -1812 1099 -1732
rect 1381 -1765 1382 -1685
rect 1384 -1765 1385 -1685
rect 1699 -1679 1739 -1678
rect 1699 -1682 1739 -1681
rect 1799 -1690 1800 -1650
rect 1802 -1690 1803 -1650
rect 1430 -1762 1431 -1722
rect 1433 -1762 1434 -1722
rect 2011 -1708 2012 -1668
rect 2014 -1708 2015 -1668
rect 2063 -1708 2064 -1668
rect 2066 -1708 2067 -1668
rect 1699 -1730 1739 -1729
rect 1699 -1733 1739 -1732
rect 562 -1950 563 -1910
rect 565 -1950 566 -1910
rect 589 -1950 590 -1910
rect 592 -1950 593 -1910
rect 873 -1907 874 -1867
rect 876 -1907 877 -1867
rect 1095 -1912 1096 -1832
rect 1098 -1912 1099 -1832
rect 1144 -1909 1145 -1869
rect 1147 -1909 1148 -1869
rect 624 -2020 625 -1980
rect 627 -2020 628 -1980
rect 550 -2199 551 -2159
rect 553 -2199 554 -2159
rect 577 -2199 578 -2159
rect 580 -2199 581 -2159
rect 612 -2269 613 -2229
rect 615 -2269 616 -2229
rect -339 -2384 -338 -2344
rect -336 -2384 -335 -2344
rect -287 -2384 -286 -2344
rect -284 -2384 -283 -2344
rect -235 -2384 -234 -2344
rect -232 -2384 -231 -2344
rect -183 -2384 -182 -2344
rect -180 -2384 -179 -2344
rect -138 -2376 -137 -2336
rect -135 -2376 -134 -2336
rect -106 -2376 -105 -2336
rect -103 -2376 -102 -2336
rect -339 -2446 -338 -2406
rect -336 -2446 -335 -2406
rect -287 -2446 -286 -2406
rect -284 -2446 -283 -2406
rect 152 -2513 192 -2512
rect 152 -2516 192 -2515
rect 252 -2524 253 -2484
rect 255 -2524 256 -2484
rect 643 -2546 644 -2506
rect 646 -2546 647 -2506
rect 670 -2546 671 -2506
rect 673 -2546 674 -2506
rect 152 -2564 192 -2563
rect 152 -2567 192 -2566
rect -339 -2654 -338 -2614
rect -336 -2654 -335 -2614
rect -287 -2654 -286 -2614
rect -284 -2654 -283 -2614
rect -235 -2654 -234 -2614
rect -232 -2654 -231 -2614
rect -183 -2654 -182 -2614
rect -180 -2654 -179 -2614
rect -138 -2646 -137 -2606
rect -135 -2646 -134 -2606
rect -106 -2646 -105 -2606
rect -103 -2646 -102 -2606
rect -339 -2716 -338 -2676
rect -336 -2716 -335 -2676
rect -287 -2716 -286 -2676
rect -284 -2716 -283 -2676
rect 169 -2668 170 -2628
rect 172 -2668 173 -2628
rect 196 -2668 197 -2628
rect 199 -2668 200 -2628
rect 705 -2616 706 -2576
rect 708 -2616 709 -2576
rect 978 -2598 979 -2558
rect 981 -2598 982 -2558
rect 1005 -2598 1006 -2558
rect 1008 -2598 1009 -2558
rect 1308 -2579 1309 -2499
rect 1311 -2579 1312 -2499
rect 1040 -2668 1041 -2628
rect 1043 -2668 1044 -2628
rect 1308 -2679 1309 -2599
rect 1311 -2679 1312 -2599
rect 231 -2738 232 -2698
rect 234 -2738 235 -2698
rect 1357 -2676 1358 -2636
rect 1360 -2676 1361 -2636
rect 644 -2829 645 -2789
rect 647 -2829 648 -2789
rect 671 -2829 672 -2789
rect 674 -2829 675 -2789
rect 706 -2899 707 -2859
rect 709 -2899 710 -2859
rect 979 -2881 980 -2841
rect 982 -2881 983 -2841
rect 1006 -2881 1007 -2841
rect 1009 -2881 1010 -2841
rect 1041 -2951 1042 -2911
rect 1044 -2951 1045 -2911
rect 1315 -2968 1316 -2888
rect 1318 -2968 1319 -2888
rect 1812 -2893 1813 -2813
rect 1815 -2893 1816 -2813
rect 2085 -2888 2086 -2848
rect 2088 -2888 2089 -2848
rect 2137 -2888 2138 -2848
rect 2140 -2888 2141 -2848
rect 2189 -2888 2190 -2848
rect 2192 -2888 2193 -2848
rect 2241 -2888 2242 -2848
rect 2244 -2888 2245 -2848
rect 2286 -2880 2287 -2840
rect 2289 -2880 2290 -2840
rect 2318 -2880 2319 -2840
rect 2321 -2880 2322 -2840
rect 640 -3100 641 -3060
rect 643 -3100 644 -3060
rect 667 -3100 668 -3060
rect 670 -3100 671 -3060
rect 1315 -3068 1316 -2988
rect 1318 -3068 1319 -2988
rect 1812 -2993 1813 -2913
rect 1815 -2993 1816 -2913
rect 2085 -2950 2086 -2910
rect 2088 -2950 2089 -2910
rect 2137 -2950 2138 -2910
rect 2140 -2950 2141 -2910
rect 1861 -2990 1862 -2950
rect 1864 -2990 1865 -2950
rect 1364 -3065 1365 -3025
rect 1367 -3065 1368 -3025
rect 1607 -3124 1608 -3044
rect 1610 -3124 1611 -3044
rect 702 -3170 703 -3130
rect 705 -3170 706 -3130
rect 1607 -3224 1608 -3144
rect 1610 -3224 1611 -3144
rect 1309 -3283 1310 -3243
rect 1312 -3283 1313 -3243
rect 1336 -3283 1337 -3243
rect 1339 -3283 1340 -3243
rect 1656 -3221 1657 -3181
rect 1659 -3221 1660 -3181
rect 628 -3349 629 -3309
rect 631 -3349 632 -3309
rect 655 -3349 656 -3309
rect 658 -3349 659 -3309
rect 1371 -3353 1372 -3313
rect 1374 -3353 1375 -3313
rect 690 -3419 691 -3379
rect 693 -3419 694 -3379
rect 969 -3415 970 -3375
rect 972 -3415 973 -3375
rect 996 -3415 997 -3375
rect 999 -3415 1000 -3375
rect 1031 -3485 1032 -3445
rect 1034 -3485 1035 -3445
rect 645 -3616 646 -3576
rect 648 -3616 649 -3576
rect 672 -3616 673 -3576
rect 675 -3616 676 -3576
rect 707 -3686 708 -3646
rect 710 -3686 711 -3646
rect 633 -3865 634 -3825
rect 636 -3865 637 -3825
rect 660 -3865 661 -3825
rect 663 -3865 664 -3825
rect 695 -3935 696 -3895
rect 698 -3935 699 -3895
<< ndcontact >>
rect 774 1646 794 1650
rect 774 1638 794 1642
rect 872 1631 876 1651
rect 880 1631 884 1651
rect 774 1595 794 1599
rect 872 1598 876 1618
rect 880 1598 884 1618
rect 908 1596 912 1616
rect 916 1596 920 1616
rect 774 1587 794 1591
rect 999 1580 1003 1600
rect 1007 1580 1011 1600
rect 1192 1575 1196 1615
rect 1200 1575 1204 1615
rect 2822 1619 2842 1623
rect 2822 1611 2842 1615
rect 2920 1604 2924 1624
rect 2928 1604 2932 1624
rect 2822 1568 2842 1572
rect 2920 1571 2924 1591
rect 2928 1571 2932 1591
rect 2956 1569 2960 1589
rect 2964 1569 2968 1589
rect 1192 1510 1196 1550
rect 1200 1510 1204 1550
rect 1235 1541 1239 1561
rect 1243 1541 1247 1561
rect 2822 1560 2842 1564
rect 3047 1553 3051 1573
rect 3055 1553 3059 1573
rect 1049 1476 1053 1496
rect 1057 1476 1061 1496
rect 1082 1476 1086 1496
rect 1090 1476 1094 1496
rect 1113 1486 1117 1506
rect 1121 1486 1125 1506
rect 3240 1548 3244 1588
rect 3248 1548 3252 1588
rect 3240 1483 3244 1523
rect 3248 1483 3252 1523
rect 3283 1514 3287 1534
rect 3291 1514 3295 1534
rect 3097 1449 3101 1469
rect 3105 1449 3109 1469
rect 3130 1449 3134 1469
rect 3138 1449 3142 1469
rect 3161 1459 3165 1479
rect 3169 1459 3173 1479
rect -1327 327 -1323 347
rect -1319 327 -1315 347
rect -1295 327 -1291 347
rect -1287 327 -1283 347
rect -1424 303 -1420 323
rect -1416 303 -1412 323
rect -1372 303 -1368 323
rect -1364 303 -1360 323
rect 3968 324 3972 344
rect 3976 324 3980 344
rect 4000 324 4004 344
rect 4008 324 4012 344
rect 3871 300 3875 320
rect 3879 300 3883 320
rect 3923 300 3927 320
rect 3931 300 3935 320
rect -1528 256 -1524 276
rect -1520 256 -1516 276
rect -1476 256 -1472 276
rect -1468 256 -1464 276
rect -1424 256 -1420 276
rect -1416 256 -1412 276
rect -1372 256 -1368 276
rect -1364 256 -1360 276
rect 3767 253 3771 273
rect 3775 253 3779 273
rect 3819 253 3823 273
rect 3827 253 3831 273
rect 3871 253 3875 273
rect 3879 253 3883 273
rect 3923 253 3927 273
rect 3931 253 3935 273
rect 1033 8 1053 12
rect 1033 0 1053 4
rect 1131 -7 1135 13
rect 1139 -7 1143 13
rect 1033 -43 1053 -39
rect 1131 -40 1135 -20
rect 1139 -40 1143 -20
rect 1620 21 1624 41
rect 1628 21 1632 41
rect 1652 21 1656 41
rect 1660 21 1664 41
rect 1523 -3 1527 17
rect 1531 -3 1535 17
rect 1575 -3 1579 17
rect 1583 -3 1587 17
rect 1167 -42 1171 -22
rect 1175 -42 1179 -22
rect 1033 -51 1053 -47
rect -201 -74 -197 -54
rect -193 -74 -189 -54
rect -169 -74 -165 -54
rect -161 -74 -157 -54
rect 1419 -50 1423 -30
rect 1427 -50 1431 -30
rect 1471 -50 1475 -30
rect 1479 -50 1483 -30
rect 1523 -50 1527 -30
rect 1531 -50 1535 -30
rect 1575 -50 1579 -30
rect 1583 -50 1587 -30
rect -298 -98 -294 -78
rect -290 -98 -286 -78
rect -246 -98 -242 -78
rect -238 -98 -234 -78
rect -402 -145 -398 -125
rect -394 -145 -390 -125
rect -350 -145 -346 -125
rect -342 -145 -338 -125
rect -298 -145 -294 -125
rect -290 -145 -286 -125
rect -246 -145 -242 -125
rect -238 -145 -234 -125
rect 120 -191 140 -187
rect 120 -199 140 -195
rect 218 -206 222 -186
rect 226 -206 230 -186
rect 120 -242 140 -238
rect 218 -239 222 -219
rect 226 -239 230 -219
rect 254 -241 258 -221
rect 262 -241 266 -221
rect 120 -250 140 -246
rect 465 -259 469 -219
rect 473 -259 477 -219
rect 1028 -212 1048 -208
rect 1028 -220 1048 -216
rect 1126 -227 1130 -207
rect 1134 -227 1138 -207
rect -205 -329 -201 -309
rect -197 -329 -193 -309
rect -173 -329 -169 -309
rect -165 -329 -161 -309
rect -302 -353 -298 -333
rect -294 -353 -290 -333
rect -250 -353 -246 -333
rect -242 -353 -238 -333
rect 465 -324 469 -284
rect 473 -324 477 -284
rect 508 -293 512 -273
rect 516 -293 520 -273
rect 801 -285 805 -265
rect 809 -285 813 -265
rect 834 -285 838 -265
rect 842 -285 846 -265
rect 865 -275 869 -255
rect 873 -275 877 -255
rect 1028 -263 1048 -259
rect 1126 -260 1130 -240
rect 1134 -260 1138 -240
rect 1162 -262 1166 -242
rect 1170 -262 1174 -242
rect 1028 -271 1048 -267
rect 1635 -255 1639 -235
rect 1643 -255 1647 -235
rect 1667 -255 1671 -235
rect 1675 -255 1679 -235
rect 1538 -279 1542 -259
rect 1546 -279 1550 -259
rect 1590 -279 1594 -259
rect 1598 -279 1602 -259
rect 1434 -326 1438 -306
rect 1442 -326 1446 -306
rect 1486 -326 1490 -306
rect 1494 -326 1498 -306
rect 1538 -326 1542 -306
rect 1546 -326 1550 -306
rect 1590 -326 1594 -306
rect 1598 -326 1602 -306
rect -406 -400 -402 -380
rect -398 -400 -394 -380
rect -354 -400 -350 -380
rect -346 -400 -342 -380
rect -302 -400 -298 -380
rect -294 -400 -290 -380
rect -250 -400 -246 -380
rect -242 -400 -238 -380
rect 190 -421 194 -381
rect 198 -421 202 -381
rect 190 -486 194 -446
rect 198 -486 202 -446
rect 233 -455 237 -435
rect 241 -455 245 -435
rect -108 -911 -104 -891
rect -100 -911 -96 -891
rect -76 -911 -72 -891
rect -68 -911 -64 -891
rect 645 -910 649 -870
rect 653 -910 657 -870
rect -205 -935 -201 -915
rect -197 -935 -193 -915
rect -153 -935 -149 -915
rect -145 -935 -141 -915
rect -309 -982 -305 -962
rect -301 -982 -297 -962
rect -257 -982 -253 -962
rect -249 -982 -245 -962
rect -205 -982 -201 -962
rect -197 -982 -193 -962
rect -153 -982 -149 -962
rect -145 -982 -141 -962
rect 108 -977 128 -973
rect 108 -985 128 -981
rect 206 -992 210 -972
rect 214 -992 218 -972
rect 645 -975 649 -935
rect 653 -975 657 -935
rect 688 -944 692 -924
rect 696 -944 700 -924
rect 945 -932 949 -912
rect 953 -932 957 -912
rect 978 -932 982 -912
rect 986 -932 990 -912
rect 1009 -922 1013 -902
rect 1017 -922 1021 -902
rect 1196 -934 1200 -914
rect 1204 -934 1208 -914
rect 1229 -934 1233 -914
rect 1237 -934 1241 -914
rect 1260 -924 1264 -904
rect 1268 -924 1272 -904
rect 1480 -942 1500 -938
rect 1480 -950 1500 -946
rect 1578 -957 1582 -937
rect 1586 -957 1590 -937
rect 108 -1028 128 -1024
rect 206 -1025 210 -1005
rect 214 -1025 218 -1005
rect 1480 -993 1500 -989
rect 1578 -990 1582 -970
rect 1586 -990 1590 -970
rect 2019 -928 2023 -908
rect 2027 -928 2031 -908
rect 2051 -928 2055 -908
rect 2059 -928 2063 -908
rect 1922 -952 1926 -932
rect 1930 -952 1934 -932
rect 1974 -952 1978 -932
rect 1982 -952 1986 -932
rect 1614 -992 1618 -972
rect 1622 -992 1626 -972
rect 1480 -1001 1500 -997
rect 1818 -999 1822 -979
rect 1826 -999 1830 -979
rect 1870 -999 1874 -979
rect 1878 -999 1882 -979
rect 1922 -999 1926 -979
rect 1930 -999 1934 -979
rect 1974 -999 1978 -979
rect 1982 -999 1986 -979
rect 242 -1027 246 -1007
rect 250 -1027 254 -1007
rect 108 -1036 128 -1032
rect -3579 -1211 -3559 -1207
rect -3579 -1219 -3559 -1215
rect -3481 -1226 -3477 -1206
rect -3473 -1226 -3469 -1206
rect -3579 -1262 -3559 -1258
rect -3481 -1259 -3477 -1239
rect -3473 -1259 -3469 -1239
rect -127 -1134 -123 -1114
rect -119 -1134 -115 -1114
rect -95 -1134 -91 -1114
rect -87 -1134 -83 -1114
rect -224 -1158 -220 -1138
rect -216 -1158 -212 -1138
rect -172 -1158 -168 -1138
rect -164 -1158 -160 -1138
rect -328 -1205 -324 -1185
rect -320 -1205 -316 -1185
rect -276 -1205 -272 -1185
rect -268 -1205 -264 -1185
rect -224 -1205 -220 -1185
rect -216 -1205 -212 -1185
rect -172 -1205 -168 -1185
rect -164 -1205 -160 -1185
rect -3445 -1261 -3441 -1241
rect -3437 -1261 -3433 -1241
rect 178 -1207 182 -1167
rect 186 -1207 190 -1167
rect -3579 -1270 -3559 -1266
rect -3354 -1277 -3350 -1257
rect -3346 -1277 -3342 -1257
rect -3161 -1282 -3157 -1242
rect -3153 -1282 -3149 -1242
rect 568 -1155 572 -1115
rect 576 -1155 580 -1115
rect 786 -1155 790 -1115
rect 794 -1155 798 -1115
rect 568 -1220 572 -1180
rect 576 -1220 580 -1180
rect 611 -1189 615 -1169
rect 619 -1189 623 -1169
rect 786 -1220 790 -1180
rect 794 -1220 798 -1180
rect 829 -1189 833 -1169
rect 837 -1189 841 -1169
rect 178 -1272 182 -1232
rect 186 -1272 190 -1232
rect 221 -1241 225 -1221
rect 229 -1241 233 -1221
rect -3161 -1347 -3157 -1307
rect -3153 -1347 -3149 -1307
rect -3118 -1316 -3114 -1296
rect -3110 -1316 -3106 -1296
rect -3304 -1381 -3300 -1361
rect -3296 -1381 -3292 -1361
rect -3271 -1381 -3267 -1361
rect -3263 -1381 -3259 -1361
rect -3240 -1371 -3236 -1351
rect -3232 -1371 -3228 -1351
rect -127 -1472 -123 -1452
rect -119 -1472 -115 -1452
rect -95 -1472 -91 -1452
rect -87 -1472 -83 -1452
rect 580 -1470 584 -1430
rect 588 -1470 592 -1430
rect -224 -1496 -220 -1476
rect -216 -1496 -212 -1476
rect -172 -1496 -168 -1476
rect -164 -1496 -160 -1476
rect -328 -1543 -324 -1523
rect -320 -1543 -316 -1523
rect -276 -1543 -272 -1523
rect -268 -1543 -264 -1523
rect -224 -1543 -220 -1523
rect -216 -1543 -212 -1523
rect -172 -1543 -168 -1523
rect -164 -1543 -160 -1523
rect 580 -1535 584 -1495
rect 588 -1535 592 -1495
rect 623 -1504 627 -1484
rect 631 -1504 635 -1484
rect 117 -1637 137 -1633
rect 117 -1645 137 -1641
rect 215 -1652 219 -1632
rect 223 -1652 227 -1632
rect 117 -1688 137 -1684
rect 215 -1685 219 -1665
rect 223 -1685 227 -1665
rect 251 -1687 255 -1667
rect 259 -1687 263 -1667
rect 117 -1696 137 -1692
rect 581 -1753 585 -1713
rect 589 -1753 593 -1713
rect -142 -1809 -138 -1789
rect -134 -1809 -130 -1789
rect -110 -1809 -106 -1789
rect -102 -1809 -98 -1789
rect 817 -1700 821 -1660
rect 825 -1700 829 -1660
rect 1065 -1657 1069 -1637
rect 1073 -1657 1077 -1637
rect 1098 -1657 1102 -1637
rect 1106 -1657 1110 -1637
rect 1129 -1647 1133 -1627
rect 1137 -1647 1141 -1627
rect 817 -1765 821 -1725
rect 825 -1765 829 -1725
rect 860 -1734 864 -1714
rect 868 -1734 872 -1714
rect -239 -1833 -235 -1813
rect -231 -1833 -227 -1813
rect -187 -1833 -183 -1813
rect -179 -1833 -175 -1813
rect -343 -1880 -339 -1860
rect -335 -1880 -331 -1860
rect -291 -1880 -287 -1860
rect -283 -1880 -279 -1860
rect -239 -1880 -235 -1860
rect -231 -1880 -227 -1860
rect -187 -1880 -183 -1860
rect -179 -1880 -175 -1860
rect 187 -1867 191 -1827
rect 195 -1867 199 -1827
rect 581 -1818 585 -1778
rect 589 -1818 593 -1778
rect 624 -1787 628 -1767
rect 632 -1787 636 -1767
rect 1661 -1678 1681 -1674
rect 1661 -1686 1681 -1682
rect 1759 -1693 1763 -1673
rect 1767 -1693 1771 -1673
rect 1661 -1729 1681 -1725
rect 1759 -1726 1763 -1706
rect 1767 -1726 1771 -1706
rect 2208 -1678 2212 -1658
rect 2216 -1678 2220 -1658
rect 2240 -1678 2244 -1658
rect 2248 -1678 2252 -1658
rect 2111 -1702 2115 -1682
rect 2119 -1702 2123 -1682
rect 2163 -1702 2167 -1682
rect 2171 -1702 2175 -1682
rect 1795 -1728 1799 -1708
rect 1803 -1728 1807 -1708
rect 1661 -1737 1681 -1733
rect 2007 -1749 2011 -1729
rect 2015 -1749 2019 -1729
rect 2059 -1749 2063 -1729
rect 2067 -1749 2071 -1729
rect 2111 -1749 2115 -1729
rect 2119 -1749 2123 -1729
rect 2163 -1749 2167 -1729
rect 2171 -1749 2175 -1729
rect 1362 -1810 1366 -1790
rect 1370 -1810 1374 -1790
rect 1395 -1810 1399 -1790
rect 1403 -1810 1407 -1790
rect 1426 -1800 1430 -1780
rect 1434 -1800 1438 -1780
rect 187 -1932 191 -1892
rect 195 -1932 199 -1892
rect 230 -1901 234 -1881
rect 238 -1901 242 -1881
rect 826 -1911 830 -1871
rect 834 -1911 838 -1871
rect 577 -2024 581 -1984
rect 585 -2024 589 -1984
rect 826 -1976 830 -1936
rect 834 -1976 838 -1936
rect 869 -1945 873 -1925
rect 877 -1945 881 -1925
rect 1076 -1957 1080 -1937
rect 1084 -1957 1088 -1937
rect 1109 -1957 1113 -1937
rect 1117 -1957 1121 -1937
rect 1140 -1947 1144 -1927
rect 1148 -1947 1152 -1927
rect 577 -2089 581 -2049
rect 585 -2089 589 -2049
rect 620 -2058 624 -2038
rect 628 -2058 632 -2038
rect 565 -2273 569 -2233
rect 573 -2273 577 -2233
rect 565 -2338 569 -2298
rect 573 -2338 577 -2298
rect 608 -2307 612 -2287
rect 616 -2307 620 -2287
rect -142 -2416 -138 -2396
rect -134 -2416 -130 -2396
rect -110 -2416 -106 -2396
rect -102 -2416 -98 -2396
rect -239 -2440 -235 -2420
rect -231 -2440 -227 -2420
rect -187 -2440 -183 -2420
rect -179 -2440 -175 -2420
rect -343 -2487 -339 -2467
rect -335 -2487 -331 -2467
rect -291 -2487 -287 -2467
rect -283 -2487 -279 -2467
rect -239 -2487 -235 -2467
rect -231 -2487 -227 -2467
rect -187 -2487 -183 -2467
rect -179 -2487 -175 -2467
rect 114 -2512 134 -2508
rect 114 -2520 134 -2516
rect 212 -2527 216 -2507
rect 220 -2527 224 -2507
rect 114 -2563 134 -2559
rect 212 -2560 216 -2540
rect 220 -2560 224 -2540
rect 248 -2562 252 -2542
rect 256 -2562 260 -2542
rect 114 -2571 134 -2567
rect 658 -2620 662 -2580
rect 666 -2620 670 -2580
rect -142 -2686 -138 -2666
rect -134 -2686 -130 -2666
rect -110 -2686 -106 -2666
rect -102 -2686 -98 -2666
rect -239 -2710 -235 -2690
rect -231 -2710 -227 -2690
rect -187 -2710 -183 -2690
rect -179 -2710 -175 -2690
rect -343 -2757 -339 -2737
rect -335 -2757 -331 -2737
rect -291 -2757 -287 -2737
rect -283 -2757 -279 -2737
rect -239 -2757 -235 -2737
rect -231 -2757 -227 -2737
rect -187 -2757 -183 -2737
rect -179 -2757 -175 -2737
rect 184 -2742 188 -2702
rect 192 -2742 196 -2702
rect 658 -2685 662 -2645
rect 666 -2685 670 -2645
rect 701 -2654 705 -2634
rect 709 -2654 713 -2634
rect 993 -2672 997 -2632
rect 1001 -2672 1005 -2632
rect 993 -2737 997 -2697
rect 1001 -2737 1005 -2697
rect 1036 -2706 1040 -2686
rect 1044 -2706 1048 -2686
rect 1289 -2724 1293 -2704
rect 1297 -2724 1301 -2704
rect 1322 -2724 1326 -2704
rect 1330 -2724 1334 -2704
rect 1353 -2714 1357 -2694
rect 1361 -2714 1365 -2694
rect 184 -2807 188 -2767
rect 192 -2807 196 -2767
rect 227 -2776 231 -2756
rect 235 -2776 239 -2756
rect 659 -2903 663 -2863
rect 667 -2903 671 -2863
rect 659 -2968 663 -2928
rect 667 -2968 671 -2928
rect 702 -2937 706 -2917
rect 710 -2937 714 -2917
rect 994 -2955 998 -2915
rect 1002 -2955 1006 -2915
rect 994 -3020 998 -2980
rect 1002 -3020 1006 -2980
rect 1037 -2989 1041 -2969
rect 1045 -2989 1049 -2969
rect 2282 -2920 2286 -2900
rect 2290 -2920 2294 -2900
rect 2314 -2920 2318 -2900
rect 2322 -2920 2326 -2900
rect 2185 -2944 2189 -2924
rect 2193 -2944 2197 -2924
rect 2237 -2944 2241 -2924
rect 2245 -2944 2249 -2924
rect 2081 -2991 2085 -2971
rect 2089 -2991 2093 -2971
rect 2133 -2991 2137 -2971
rect 2141 -2991 2145 -2971
rect 2185 -2991 2189 -2971
rect 2193 -2991 2197 -2971
rect 2237 -2991 2241 -2971
rect 2245 -2991 2249 -2971
rect 1793 -3038 1797 -3018
rect 1801 -3038 1805 -3018
rect 1826 -3038 1830 -3018
rect 1834 -3038 1838 -3018
rect 1857 -3028 1861 -3008
rect 1865 -3028 1869 -3008
rect 1296 -3113 1300 -3093
rect 1304 -3113 1308 -3093
rect 1329 -3113 1333 -3093
rect 1337 -3113 1341 -3093
rect 1360 -3103 1364 -3083
rect 1368 -3103 1372 -3083
rect 655 -3174 659 -3134
rect 663 -3174 667 -3134
rect 655 -3239 659 -3199
rect 663 -3239 667 -3199
rect 698 -3208 702 -3188
rect 706 -3208 710 -3188
rect 1588 -3269 1592 -3249
rect 1596 -3269 1600 -3249
rect 1621 -3269 1625 -3249
rect 1629 -3269 1633 -3249
rect 1652 -3259 1656 -3239
rect 1660 -3259 1664 -3239
rect 1324 -3357 1328 -3317
rect 1332 -3357 1336 -3317
rect 643 -3423 647 -3383
rect 651 -3423 655 -3383
rect 643 -3488 647 -3448
rect 651 -3488 655 -3448
rect 686 -3457 690 -3437
rect 694 -3457 698 -3437
rect 1324 -3422 1328 -3382
rect 1332 -3422 1336 -3382
rect 1367 -3391 1371 -3371
rect 1375 -3391 1379 -3371
rect 984 -3489 988 -3449
rect 992 -3489 996 -3449
rect 984 -3554 988 -3514
rect 992 -3554 996 -3514
rect 1027 -3523 1031 -3503
rect 1035 -3523 1039 -3503
rect 660 -3690 664 -3650
rect 668 -3690 672 -3650
rect 660 -3755 664 -3715
rect 668 -3755 672 -3715
rect 703 -3724 707 -3704
rect 711 -3724 715 -3704
rect 648 -3939 652 -3899
rect 656 -3939 660 -3899
rect 648 -4004 652 -3964
rect 656 -4004 660 -3964
rect 691 -3973 695 -3953
rect 699 -3973 703 -3953
<< pdcontact >>
rect 812 1646 852 1650
rect 812 1638 852 1642
rect 908 1634 912 1674
rect 916 1634 920 1674
rect 812 1595 852 1599
rect 999 1618 1003 1658
rect 1007 1618 1011 1658
rect 1064 1621 1068 1701
rect 1072 1621 1076 1701
rect 1173 1649 1177 1689
rect 1181 1649 1185 1689
rect 1200 1649 1204 1689
rect 1208 1649 1212 1689
rect 812 1587 852 1591
rect 1064 1521 1068 1601
rect 1072 1521 1076 1601
rect 1113 1524 1117 1564
rect 1121 1524 1125 1564
rect 1235 1579 1239 1619
rect 1243 1579 1247 1619
rect 2860 1619 2900 1623
rect 2860 1611 2900 1615
rect 2956 1607 2960 1647
rect 2964 1607 2968 1647
rect 2860 1568 2900 1572
rect 3047 1591 3051 1631
rect 3055 1591 3059 1631
rect 3112 1594 3116 1674
rect 3120 1594 3124 1674
rect 3221 1622 3225 1662
rect 3229 1622 3233 1662
rect 3248 1622 3252 1662
rect 3256 1622 3260 1662
rect 2860 1560 2900 1564
rect 3112 1494 3116 1574
rect 3120 1494 3124 1574
rect 3161 1497 3165 1537
rect 3169 1497 3173 1537
rect 3283 1552 3287 1592
rect 3291 1552 3295 1592
rect -1528 359 -1524 399
rect -1520 359 -1516 399
rect -1476 359 -1472 399
rect -1468 359 -1464 399
rect -1424 359 -1420 399
rect -1416 359 -1412 399
rect -1372 359 -1368 399
rect -1364 359 -1360 399
rect -1327 367 -1323 407
rect -1319 367 -1315 407
rect -1295 367 -1291 407
rect -1287 367 -1283 407
rect 3767 356 3771 396
rect 3775 356 3779 396
rect 3819 356 3823 396
rect 3827 356 3831 396
rect 3871 356 3875 396
rect 3879 356 3883 396
rect 3923 356 3927 396
rect 3931 356 3935 396
rect 3968 364 3972 404
rect 3976 364 3980 404
rect 4000 364 4004 404
rect 4008 364 4012 404
rect -1528 297 -1524 337
rect -1520 297 -1516 337
rect -1476 297 -1472 337
rect -1468 297 -1464 337
rect 3767 294 3771 334
rect 3775 294 3779 334
rect 3819 294 3823 334
rect 3827 294 3831 334
rect 1419 53 1423 93
rect 1427 53 1431 93
rect 1471 53 1475 93
rect 1479 53 1483 93
rect 1523 53 1527 93
rect 1531 53 1535 93
rect 1575 53 1579 93
rect 1583 53 1587 93
rect 1620 61 1624 101
rect 1628 61 1632 101
rect 1652 61 1656 101
rect 1660 61 1664 101
rect 1071 8 1111 12
rect -402 -42 -398 -2
rect -394 -42 -390 -2
rect -350 -42 -346 -2
rect -342 -42 -338 -2
rect -298 -42 -294 -2
rect -290 -42 -286 -2
rect -246 -42 -242 -2
rect -238 -42 -234 -2
rect -201 -34 -197 6
rect -193 -34 -189 6
rect -169 -34 -165 6
rect -161 -34 -157 6
rect 1071 0 1111 4
rect 1167 -4 1171 36
rect 1175 -4 1179 36
rect 1071 -43 1111 -39
rect 1419 -9 1423 31
rect 1427 -9 1431 31
rect 1471 -9 1475 31
rect 1479 -9 1483 31
rect 1071 -51 1111 -47
rect -402 -104 -398 -64
rect -394 -104 -390 -64
rect -350 -104 -346 -64
rect -342 -104 -338 -64
rect 816 -140 820 -60
rect 824 -140 828 -60
rect 158 -191 198 -187
rect 158 -199 198 -195
rect 254 -203 258 -163
rect 262 -203 266 -163
rect 446 -185 450 -145
rect 454 -185 458 -145
rect 473 -185 477 -145
rect 481 -185 485 -145
rect 158 -242 198 -238
rect -406 -297 -402 -257
rect -398 -297 -394 -257
rect -354 -297 -350 -257
rect -346 -297 -342 -257
rect -302 -297 -298 -257
rect -294 -297 -290 -257
rect -250 -297 -246 -257
rect -242 -297 -238 -257
rect -205 -289 -201 -249
rect -197 -289 -193 -249
rect -173 -289 -169 -249
rect -165 -289 -161 -249
rect 158 -250 198 -246
rect 508 -255 512 -215
rect 516 -255 520 -215
rect 816 -240 820 -160
rect 824 -240 828 -160
rect 865 -237 869 -197
rect 873 -237 877 -197
rect 1066 -212 1106 -208
rect 1066 -220 1106 -216
rect 1162 -224 1166 -184
rect 1170 -224 1174 -184
rect 1434 -223 1438 -183
rect 1442 -223 1446 -183
rect 1486 -223 1490 -183
rect 1494 -223 1498 -183
rect 1538 -223 1542 -183
rect 1546 -223 1550 -183
rect 1590 -223 1594 -183
rect 1598 -223 1602 -183
rect 1635 -215 1639 -175
rect 1643 -215 1647 -175
rect 1667 -215 1671 -175
rect 1675 -215 1679 -175
rect -406 -359 -402 -319
rect -398 -359 -394 -319
rect -354 -359 -350 -319
rect -346 -359 -342 -319
rect 171 -347 175 -307
rect 179 -347 183 -307
rect 198 -347 202 -307
rect 206 -347 210 -307
rect 1066 -263 1106 -259
rect 1066 -271 1106 -267
rect 1434 -285 1438 -245
rect 1442 -285 1446 -245
rect 1486 -285 1490 -245
rect 1494 -285 1498 -245
rect 233 -417 237 -377
rect 241 -417 245 -377
rect 960 -787 964 -707
rect 968 -787 972 -707
rect 1211 -789 1215 -709
rect 1219 -789 1223 -709
rect -309 -879 -305 -839
rect -301 -879 -297 -839
rect -257 -879 -253 -839
rect -249 -879 -245 -839
rect -205 -879 -201 -839
rect -197 -879 -193 -839
rect -153 -879 -149 -839
rect -145 -879 -141 -839
rect -108 -871 -104 -831
rect -100 -871 -96 -831
rect -76 -871 -72 -831
rect -68 -871 -64 -831
rect 626 -836 630 -796
rect 634 -836 638 -796
rect 653 -836 657 -796
rect 661 -836 665 -796
rect -309 -941 -305 -901
rect -301 -941 -297 -901
rect -257 -941 -253 -901
rect -249 -941 -245 -901
rect 688 -906 692 -866
rect 696 -906 700 -866
rect 960 -887 964 -807
rect 968 -887 972 -807
rect 1009 -884 1013 -844
rect 1017 -884 1021 -844
rect 1211 -889 1215 -809
rect 1219 -889 1223 -809
rect 146 -977 186 -973
rect 146 -985 186 -981
rect 242 -989 246 -949
rect 250 -989 254 -949
rect 1260 -886 1264 -846
rect 1268 -886 1272 -846
rect 1818 -896 1822 -856
rect 1826 -896 1830 -856
rect 1870 -896 1874 -856
rect 1878 -896 1882 -856
rect 1922 -896 1926 -856
rect 1930 -896 1934 -856
rect 1974 -896 1978 -856
rect 1982 -896 1986 -856
rect 2019 -888 2023 -848
rect 2027 -888 2031 -848
rect 2051 -888 2055 -848
rect 2059 -888 2063 -848
rect 1518 -942 1558 -938
rect 1518 -950 1558 -946
rect 1614 -954 1618 -914
rect 1622 -954 1626 -914
rect 146 -1028 186 -1024
rect 1518 -993 1558 -989
rect 1818 -958 1822 -918
rect 1826 -958 1830 -918
rect 1870 -958 1874 -918
rect 1878 -958 1882 -918
rect 1518 -1001 1558 -997
rect 146 -1036 186 -1032
rect -328 -1102 -324 -1062
rect -320 -1102 -316 -1062
rect -276 -1102 -272 -1062
rect -268 -1102 -264 -1062
rect -224 -1102 -220 -1062
rect -216 -1102 -212 -1062
rect -172 -1102 -168 -1062
rect -164 -1102 -160 -1062
rect -127 -1094 -123 -1054
rect -119 -1094 -115 -1054
rect -95 -1094 -91 -1054
rect -87 -1094 -83 -1054
rect 549 -1081 553 -1041
rect 557 -1081 561 -1041
rect 576 -1081 580 -1041
rect 584 -1081 588 -1041
rect 767 -1081 771 -1041
rect 775 -1081 779 -1041
rect 794 -1081 798 -1041
rect 802 -1081 806 -1041
rect -3541 -1211 -3501 -1207
rect -3541 -1219 -3501 -1215
rect -3445 -1223 -3441 -1183
rect -3437 -1223 -3433 -1183
rect -3541 -1262 -3501 -1258
rect -3354 -1239 -3350 -1199
rect -3346 -1239 -3342 -1199
rect -3289 -1236 -3285 -1156
rect -3281 -1236 -3277 -1156
rect -328 -1164 -324 -1124
rect -320 -1164 -316 -1124
rect -276 -1164 -272 -1124
rect -268 -1164 -264 -1124
rect 159 -1133 163 -1093
rect 167 -1133 171 -1093
rect 186 -1133 190 -1093
rect 194 -1133 198 -1093
rect -3180 -1208 -3176 -1168
rect -3172 -1208 -3168 -1168
rect -3153 -1208 -3149 -1168
rect -3145 -1208 -3141 -1168
rect -3541 -1270 -3501 -1266
rect -3289 -1336 -3285 -1256
rect -3281 -1336 -3277 -1256
rect -3240 -1333 -3236 -1293
rect -3232 -1333 -3228 -1293
rect 221 -1203 225 -1163
rect 229 -1203 233 -1163
rect 611 -1151 615 -1111
rect 619 -1151 623 -1111
rect 829 -1151 833 -1111
rect 837 -1151 841 -1111
rect -3118 -1278 -3114 -1238
rect -3110 -1278 -3106 -1238
rect -328 -1440 -324 -1400
rect -320 -1440 -316 -1400
rect -276 -1440 -272 -1400
rect -268 -1440 -264 -1400
rect -224 -1440 -220 -1400
rect -216 -1440 -212 -1400
rect -172 -1440 -168 -1400
rect -164 -1440 -160 -1400
rect -127 -1432 -123 -1392
rect -119 -1432 -115 -1392
rect -95 -1432 -91 -1392
rect -87 -1432 -83 -1392
rect 561 -1396 565 -1356
rect 569 -1396 573 -1356
rect 588 -1396 592 -1356
rect 596 -1396 600 -1356
rect -328 -1502 -324 -1462
rect -320 -1502 -316 -1462
rect -276 -1502 -272 -1462
rect -268 -1502 -264 -1462
rect 623 -1466 627 -1426
rect 631 -1466 635 -1426
rect 1080 -1512 1084 -1432
rect 1088 -1512 1092 -1432
rect 155 -1637 195 -1633
rect 155 -1645 195 -1641
rect 251 -1649 255 -1609
rect 259 -1649 263 -1609
rect 798 -1626 802 -1586
rect 806 -1626 810 -1586
rect 825 -1626 829 -1586
rect 833 -1626 837 -1586
rect 1080 -1612 1084 -1532
rect 1088 -1612 1092 -1532
rect 155 -1688 195 -1684
rect 562 -1679 566 -1639
rect 570 -1679 574 -1639
rect 589 -1679 593 -1639
rect 597 -1679 601 -1639
rect 1129 -1609 1133 -1569
rect 1137 -1609 1141 -1569
rect 155 -1696 195 -1692
rect -343 -1777 -339 -1737
rect -335 -1777 -331 -1737
rect -291 -1777 -287 -1737
rect -283 -1777 -279 -1737
rect -239 -1777 -235 -1737
rect -231 -1777 -227 -1737
rect -187 -1777 -183 -1737
rect -179 -1777 -175 -1737
rect -142 -1769 -138 -1729
rect -134 -1769 -130 -1729
rect -110 -1769 -106 -1729
rect -102 -1769 -98 -1729
rect -343 -1839 -339 -1799
rect -335 -1839 -331 -1799
rect -291 -1839 -287 -1799
rect -283 -1839 -279 -1799
rect 168 -1793 172 -1753
rect 176 -1793 180 -1753
rect 195 -1793 199 -1753
rect 203 -1793 207 -1753
rect 624 -1749 628 -1709
rect 632 -1749 636 -1709
rect 860 -1696 864 -1656
rect 868 -1696 872 -1656
rect 1377 -1665 1381 -1585
rect 1385 -1665 1389 -1585
rect 2007 -1646 2011 -1606
rect 2015 -1646 2019 -1606
rect 2059 -1646 2063 -1606
rect 2067 -1646 2071 -1606
rect 2111 -1646 2115 -1606
rect 2119 -1646 2123 -1606
rect 2163 -1646 2167 -1606
rect 2171 -1646 2175 -1606
rect 2208 -1638 2212 -1598
rect 2216 -1638 2220 -1598
rect 2240 -1638 2244 -1598
rect 2248 -1638 2252 -1598
rect 230 -1863 234 -1823
rect 238 -1863 242 -1823
rect 807 -1837 811 -1797
rect 815 -1837 819 -1797
rect 834 -1837 838 -1797
rect 842 -1837 846 -1797
rect 1091 -1812 1095 -1732
rect 1099 -1812 1103 -1732
rect 1377 -1765 1381 -1685
rect 1385 -1765 1389 -1685
rect 1699 -1678 1739 -1674
rect 1699 -1686 1739 -1682
rect 1795 -1690 1799 -1650
rect 1803 -1690 1807 -1650
rect 1426 -1762 1430 -1722
rect 1434 -1762 1438 -1722
rect 1699 -1729 1739 -1725
rect 2007 -1708 2011 -1668
rect 2015 -1708 2019 -1668
rect 2059 -1708 2063 -1668
rect 2067 -1708 2071 -1668
rect 1699 -1737 1739 -1733
rect 558 -1950 562 -1910
rect 566 -1950 570 -1910
rect 585 -1950 589 -1910
rect 593 -1950 597 -1910
rect 869 -1907 873 -1867
rect 877 -1907 881 -1867
rect 1091 -1912 1095 -1832
rect 1099 -1912 1103 -1832
rect 1140 -1909 1144 -1869
rect 1148 -1909 1152 -1869
rect 620 -2020 624 -1980
rect 628 -2020 632 -1980
rect 546 -2199 550 -2159
rect 554 -2199 558 -2159
rect 573 -2199 577 -2159
rect 581 -2199 585 -2159
rect 608 -2269 612 -2229
rect 616 -2269 620 -2229
rect -343 -2384 -339 -2344
rect -335 -2384 -331 -2344
rect -291 -2384 -287 -2344
rect -283 -2384 -279 -2344
rect -239 -2384 -235 -2344
rect -231 -2384 -227 -2344
rect -187 -2384 -183 -2344
rect -179 -2384 -175 -2344
rect -142 -2376 -138 -2336
rect -134 -2376 -130 -2336
rect -110 -2376 -106 -2336
rect -102 -2376 -98 -2336
rect -343 -2446 -339 -2406
rect -335 -2446 -331 -2406
rect -291 -2446 -287 -2406
rect -283 -2446 -279 -2406
rect 152 -2512 192 -2508
rect 152 -2520 192 -2516
rect 248 -2524 252 -2484
rect 256 -2524 260 -2484
rect 152 -2563 192 -2559
rect 639 -2546 643 -2506
rect 647 -2546 651 -2506
rect 666 -2546 670 -2506
rect 674 -2546 678 -2506
rect 152 -2571 192 -2567
rect -343 -2654 -339 -2614
rect -335 -2654 -331 -2614
rect -291 -2654 -287 -2614
rect -283 -2654 -279 -2614
rect -239 -2654 -235 -2614
rect -231 -2654 -227 -2614
rect -187 -2654 -183 -2614
rect -179 -2654 -175 -2614
rect -142 -2646 -138 -2606
rect -134 -2646 -130 -2606
rect -110 -2646 -106 -2606
rect -102 -2646 -98 -2606
rect -343 -2716 -339 -2676
rect -335 -2716 -331 -2676
rect -291 -2716 -287 -2676
rect -283 -2716 -279 -2676
rect 165 -2668 169 -2628
rect 173 -2668 177 -2628
rect 192 -2668 196 -2628
rect 200 -2668 204 -2628
rect 701 -2616 705 -2576
rect 709 -2616 713 -2576
rect 974 -2598 978 -2558
rect 982 -2598 986 -2558
rect 1001 -2598 1005 -2558
rect 1009 -2598 1013 -2558
rect 1304 -2579 1308 -2499
rect 1312 -2579 1316 -2499
rect 1036 -2668 1040 -2628
rect 1044 -2668 1048 -2628
rect 1304 -2679 1308 -2599
rect 1312 -2679 1316 -2599
rect 227 -2738 231 -2698
rect 235 -2738 239 -2698
rect 1353 -2676 1357 -2636
rect 1361 -2676 1365 -2636
rect 640 -2829 644 -2789
rect 648 -2829 652 -2789
rect 667 -2829 671 -2789
rect 675 -2829 679 -2789
rect 702 -2899 706 -2859
rect 710 -2899 714 -2859
rect 975 -2881 979 -2841
rect 983 -2881 987 -2841
rect 1002 -2881 1006 -2841
rect 1010 -2881 1014 -2841
rect 1037 -2951 1041 -2911
rect 1045 -2951 1049 -2911
rect 1311 -2968 1315 -2888
rect 1319 -2968 1323 -2888
rect 1808 -2893 1812 -2813
rect 1816 -2893 1820 -2813
rect 2081 -2888 2085 -2848
rect 2089 -2888 2093 -2848
rect 2133 -2888 2137 -2848
rect 2141 -2888 2145 -2848
rect 2185 -2888 2189 -2848
rect 2193 -2888 2197 -2848
rect 2237 -2888 2241 -2848
rect 2245 -2888 2249 -2848
rect 2282 -2880 2286 -2840
rect 2290 -2880 2294 -2840
rect 2314 -2880 2318 -2840
rect 2322 -2880 2326 -2840
rect 636 -3100 640 -3060
rect 644 -3100 648 -3060
rect 663 -3100 667 -3060
rect 671 -3100 675 -3060
rect 1311 -3068 1315 -2988
rect 1319 -3068 1323 -2988
rect 1808 -2993 1812 -2913
rect 1816 -2993 1820 -2913
rect 2081 -2950 2085 -2910
rect 2089 -2950 2093 -2910
rect 2133 -2950 2137 -2910
rect 2141 -2950 2145 -2910
rect 1857 -2990 1861 -2950
rect 1865 -2990 1869 -2950
rect 1360 -3065 1364 -3025
rect 1368 -3065 1372 -3025
rect 1603 -3124 1607 -3044
rect 1611 -3124 1615 -3044
rect 698 -3170 702 -3130
rect 706 -3170 710 -3130
rect 1603 -3224 1607 -3144
rect 1611 -3224 1615 -3144
rect 1305 -3283 1309 -3243
rect 1313 -3283 1317 -3243
rect 1332 -3283 1336 -3243
rect 1340 -3283 1344 -3243
rect 1652 -3221 1656 -3181
rect 1660 -3221 1664 -3181
rect 624 -3349 628 -3309
rect 632 -3349 636 -3309
rect 651 -3349 655 -3309
rect 659 -3349 663 -3309
rect 1367 -3353 1371 -3313
rect 1375 -3353 1379 -3313
rect 686 -3419 690 -3379
rect 694 -3419 698 -3379
rect 965 -3415 969 -3375
rect 973 -3415 977 -3375
rect 992 -3415 996 -3375
rect 1000 -3415 1004 -3375
rect 1027 -3485 1031 -3445
rect 1035 -3485 1039 -3445
rect 641 -3616 645 -3576
rect 649 -3616 653 -3576
rect 668 -3616 672 -3576
rect 676 -3616 680 -3576
rect 703 -3686 707 -3646
rect 711 -3686 715 -3646
rect 629 -3865 633 -3825
rect 637 -3865 641 -3825
rect 656 -3865 660 -3825
rect 664 -3865 668 -3825
rect 691 -3935 695 -3895
rect 699 -3935 703 -3895
<< psubstratepcontact >>
rect 763 1653 767 1657
rect 763 1632 767 1636
rect 763 1602 767 1606
rect 763 1581 767 1585
rect 901 1585 905 1589
rect 922 1585 926 1589
rect 992 1569 996 1573
rect 1013 1569 1017 1573
rect 2811 1626 2815 1630
rect 2811 1605 2815 1609
rect 2811 1575 2815 1579
rect 2811 1554 2815 1558
rect 2949 1558 2953 1562
rect 2970 1558 2974 1562
rect 3040 1542 3044 1546
rect 3061 1542 3065 1546
rect 1228 1530 1232 1534
rect 1249 1530 1253 1534
rect 1185 1499 1189 1503
rect 1206 1499 1210 1503
rect 1106 1475 1110 1479
rect 1127 1475 1131 1479
rect 3276 1503 3280 1507
rect 3297 1503 3301 1507
rect 1042 1465 1046 1469
rect 1063 1465 1067 1469
rect 1075 1465 1079 1469
rect 1096 1465 1100 1469
rect 3233 1472 3237 1476
rect 3254 1472 3258 1476
rect 3154 1448 3158 1452
rect 3175 1448 3179 1452
rect 3090 1438 3094 1442
rect 3111 1438 3115 1442
rect 3123 1438 3127 1442
rect 3144 1438 3148 1442
rect -1335 314 -1331 318
rect -1311 314 -1307 318
rect -1303 314 -1299 318
rect -1279 314 -1275 318
rect 3960 311 3964 315
rect 3984 311 3988 315
rect 3992 311 3996 315
rect 4016 311 4020 315
rect -1511 243 -1507 247
rect -1459 243 -1455 247
rect -1407 243 -1403 247
rect -1355 243 -1351 247
rect 3784 240 3788 244
rect 3836 240 3840 244
rect 3888 240 3892 244
rect 3940 240 3944 244
rect 1022 15 1026 19
rect 1022 -6 1026 -2
rect 1022 -36 1026 -32
rect 1612 8 1616 12
rect 1636 8 1640 12
rect 1644 8 1648 12
rect 1668 8 1672 12
rect 1022 -57 1026 -53
rect 1160 -53 1164 -49
rect 1181 -53 1185 -49
rect -209 -87 -205 -83
rect -185 -87 -181 -83
rect -177 -87 -173 -83
rect -153 -87 -149 -83
rect 1436 -63 1440 -59
rect 1488 -63 1492 -59
rect 1540 -63 1544 -59
rect 1592 -63 1596 -59
rect -385 -158 -381 -154
rect -333 -158 -329 -154
rect -281 -158 -277 -154
rect -229 -158 -225 -154
rect 109 -184 113 -180
rect 109 -205 113 -201
rect 109 -235 113 -231
rect 109 -256 113 -252
rect 247 -252 251 -248
rect 268 -252 272 -248
rect 1017 -205 1021 -201
rect 1017 -226 1021 -222
rect -213 -342 -209 -338
rect -189 -342 -185 -338
rect -181 -342 -177 -338
rect -157 -342 -153 -338
rect 1017 -256 1021 -252
rect 1017 -277 1021 -273
rect 1155 -273 1159 -269
rect 1176 -273 1180 -269
rect 858 -286 862 -282
rect 879 -286 883 -282
rect 1627 -268 1631 -264
rect 1651 -268 1655 -264
rect 1659 -268 1663 -264
rect 1683 -268 1687 -264
rect 794 -296 798 -292
rect 815 -296 819 -292
rect 827 -296 831 -292
rect 848 -296 852 -292
rect 501 -304 505 -300
rect 522 -304 526 -300
rect 458 -335 462 -331
rect 479 -335 483 -331
rect 1451 -339 1455 -335
rect 1503 -339 1507 -335
rect 1555 -339 1559 -335
rect 1607 -339 1611 -335
rect -389 -413 -385 -409
rect -337 -413 -333 -409
rect -285 -413 -281 -409
rect -233 -413 -229 -409
rect 226 -466 230 -462
rect 247 -466 251 -462
rect 183 -497 187 -493
rect 204 -497 208 -493
rect -116 -924 -112 -920
rect -92 -924 -88 -920
rect -84 -924 -80 -920
rect -60 -924 -56 -920
rect 97 -970 101 -966
rect 97 -991 101 -987
rect -292 -995 -288 -991
rect -240 -995 -236 -991
rect -188 -995 -184 -991
rect -136 -995 -132 -991
rect 1002 -933 1006 -929
rect 1023 -933 1027 -929
rect 1253 -935 1257 -931
rect 1274 -935 1278 -931
rect 1469 -935 1473 -931
rect 938 -943 942 -939
rect 959 -943 963 -939
rect 971 -943 975 -939
rect 992 -943 996 -939
rect 1189 -945 1193 -941
rect 1210 -945 1214 -941
rect 1222 -945 1226 -941
rect 1243 -945 1247 -941
rect 681 -955 685 -951
rect 702 -955 706 -951
rect 1469 -956 1473 -952
rect 638 -986 642 -982
rect 659 -986 663 -982
rect 1469 -986 1473 -982
rect 97 -1021 101 -1017
rect 2011 -941 2015 -937
rect 2035 -941 2039 -937
rect 2043 -941 2047 -937
rect 2067 -941 2071 -937
rect 1469 -1007 1473 -1003
rect 1607 -1003 1611 -999
rect 1628 -1003 1632 -999
rect 1835 -1012 1839 -1008
rect 1887 -1012 1891 -1008
rect 1939 -1012 1943 -1008
rect 1991 -1012 1995 -1008
rect 97 -1042 101 -1038
rect 235 -1038 239 -1034
rect 256 -1038 260 -1034
rect -3590 -1204 -3586 -1200
rect -3590 -1225 -3586 -1221
rect -3590 -1255 -3586 -1251
rect -135 -1147 -131 -1143
rect -111 -1147 -107 -1143
rect -103 -1147 -99 -1143
rect -79 -1147 -75 -1143
rect -311 -1218 -307 -1214
rect -259 -1218 -255 -1214
rect -207 -1218 -203 -1214
rect -155 -1218 -151 -1214
rect -3590 -1276 -3586 -1272
rect -3452 -1272 -3448 -1268
rect -3431 -1272 -3427 -1268
rect -3361 -1288 -3357 -1284
rect -3340 -1288 -3336 -1284
rect 604 -1200 608 -1196
rect 625 -1200 629 -1196
rect 822 -1200 826 -1196
rect 843 -1200 847 -1196
rect 561 -1231 565 -1227
rect 582 -1231 586 -1227
rect 779 -1231 783 -1227
rect 800 -1231 804 -1227
rect 214 -1252 218 -1248
rect 235 -1252 239 -1248
rect 171 -1283 175 -1279
rect 192 -1283 196 -1279
rect -3125 -1327 -3121 -1323
rect -3104 -1327 -3100 -1323
rect -3168 -1358 -3164 -1354
rect -3147 -1358 -3143 -1354
rect -3247 -1382 -3243 -1378
rect -3226 -1382 -3222 -1378
rect -3311 -1392 -3307 -1388
rect -3290 -1392 -3286 -1388
rect -3278 -1392 -3274 -1388
rect -3257 -1392 -3253 -1388
rect -135 -1485 -131 -1481
rect -111 -1485 -107 -1481
rect -103 -1485 -99 -1481
rect -79 -1485 -75 -1481
rect 616 -1515 620 -1511
rect 637 -1515 641 -1511
rect 573 -1546 577 -1542
rect 594 -1546 598 -1542
rect -311 -1556 -307 -1552
rect -259 -1556 -255 -1552
rect -207 -1556 -203 -1552
rect -155 -1556 -151 -1552
rect 106 -1630 110 -1626
rect 106 -1651 110 -1647
rect 106 -1681 110 -1677
rect 106 -1702 110 -1698
rect 244 -1698 248 -1694
rect 265 -1698 269 -1694
rect 1122 -1658 1126 -1654
rect 1143 -1658 1147 -1654
rect 1058 -1668 1062 -1664
rect 1079 -1668 1083 -1664
rect 1091 -1668 1095 -1664
rect 1112 -1668 1116 -1664
rect 1650 -1671 1654 -1667
rect 853 -1745 857 -1741
rect 874 -1745 878 -1741
rect -150 -1822 -146 -1818
rect -126 -1822 -122 -1818
rect -118 -1822 -114 -1818
rect -94 -1822 -90 -1818
rect 810 -1776 814 -1772
rect 831 -1776 835 -1772
rect 617 -1798 621 -1794
rect 638 -1798 642 -1794
rect 574 -1829 578 -1825
rect 595 -1829 599 -1825
rect 1650 -1692 1654 -1688
rect 1650 -1722 1654 -1718
rect 2200 -1691 2204 -1687
rect 2224 -1691 2228 -1687
rect 2232 -1691 2236 -1687
rect 2256 -1691 2260 -1687
rect 1650 -1743 1654 -1739
rect 1788 -1739 1792 -1735
rect 1809 -1739 1813 -1735
rect 2024 -1762 2028 -1758
rect 2076 -1762 2080 -1758
rect 2128 -1762 2132 -1758
rect 2180 -1762 2184 -1758
rect 1419 -1811 1423 -1807
rect 1440 -1811 1444 -1807
rect -326 -1893 -322 -1889
rect -274 -1893 -270 -1889
rect -222 -1893 -218 -1889
rect -170 -1893 -166 -1889
rect 223 -1912 227 -1908
rect 244 -1912 248 -1908
rect 180 -1943 184 -1939
rect 201 -1943 205 -1939
rect 1355 -1821 1359 -1817
rect 1376 -1821 1380 -1817
rect 1388 -1821 1392 -1817
rect 1409 -1821 1413 -1817
rect 862 -1956 866 -1952
rect 883 -1956 887 -1952
rect 1133 -1958 1137 -1954
rect 1154 -1958 1158 -1954
rect 1069 -1968 1073 -1964
rect 1090 -1968 1094 -1964
rect 1102 -1968 1106 -1964
rect 1123 -1968 1127 -1964
rect 819 -1987 823 -1983
rect 840 -1987 844 -1983
rect 613 -2069 617 -2065
rect 634 -2069 638 -2065
rect 570 -2100 574 -2096
rect 591 -2100 595 -2096
rect 601 -2318 605 -2314
rect 622 -2318 626 -2314
rect 558 -2349 562 -2345
rect 579 -2349 583 -2345
rect -150 -2429 -146 -2425
rect -126 -2429 -122 -2425
rect -118 -2429 -114 -2425
rect -94 -2429 -90 -2425
rect -326 -2500 -322 -2496
rect -274 -2500 -270 -2496
rect -222 -2500 -218 -2496
rect -170 -2500 -166 -2496
rect 103 -2505 107 -2501
rect 103 -2526 107 -2522
rect 103 -2556 107 -2552
rect 103 -2577 107 -2573
rect 241 -2573 245 -2569
rect 262 -2573 266 -2569
rect -150 -2699 -146 -2695
rect -126 -2699 -122 -2695
rect -118 -2699 -114 -2695
rect -94 -2699 -90 -2695
rect 694 -2665 698 -2661
rect 715 -2665 719 -2661
rect 651 -2696 655 -2692
rect 672 -2696 676 -2692
rect 1029 -2717 1033 -2713
rect 1050 -2717 1054 -2713
rect 1346 -2725 1350 -2721
rect 1367 -2725 1371 -2721
rect 1282 -2735 1286 -2731
rect 1303 -2735 1307 -2731
rect 1315 -2735 1319 -2731
rect 1336 -2735 1340 -2731
rect 986 -2748 990 -2744
rect 1007 -2748 1011 -2744
rect -326 -2770 -322 -2766
rect -274 -2770 -270 -2766
rect -222 -2770 -218 -2766
rect -170 -2770 -166 -2766
rect 220 -2787 224 -2783
rect 241 -2787 245 -2783
rect 177 -2818 181 -2814
rect 198 -2818 202 -2814
rect 695 -2948 699 -2944
rect 716 -2948 720 -2944
rect 652 -2979 656 -2975
rect 673 -2979 677 -2975
rect 1030 -3000 1034 -2996
rect 1051 -3000 1055 -2996
rect 987 -3031 991 -3027
rect 1008 -3031 1012 -3027
rect 2274 -2933 2278 -2929
rect 2298 -2933 2302 -2929
rect 2306 -2933 2310 -2929
rect 2330 -2933 2334 -2929
rect 2098 -3004 2102 -3000
rect 2150 -3004 2154 -3000
rect 2202 -3004 2206 -3000
rect 2254 -3004 2258 -3000
rect 1850 -3039 1854 -3035
rect 1871 -3039 1875 -3035
rect 1353 -3114 1357 -3110
rect 1374 -3114 1378 -3110
rect 1289 -3124 1293 -3120
rect 1310 -3124 1314 -3120
rect 1322 -3124 1326 -3120
rect 1343 -3124 1347 -3120
rect 1786 -3049 1790 -3045
rect 1807 -3049 1811 -3045
rect 1819 -3049 1823 -3045
rect 1840 -3049 1844 -3045
rect 691 -3219 695 -3215
rect 712 -3219 716 -3215
rect 648 -3250 652 -3246
rect 669 -3250 673 -3246
rect 1645 -3270 1649 -3266
rect 1666 -3270 1670 -3266
rect 1581 -3280 1585 -3276
rect 1602 -3280 1606 -3276
rect 1614 -3280 1618 -3276
rect 1635 -3280 1639 -3276
rect 1360 -3402 1364 -3398
rect 1381 -3402 1385 -3398
rect 679 -3468 683 -3464
rect 700 -3468 704 -3464
rect 636 -3499 640 -3495
rect 657 -3499 661 -3495
rect 1317 -3433 1321 -3429
rect 1338 -3433 1342 -3429
rect 1020 -3534 1024 -3530
rect 1041 -3534 1045 -3530
rect 977 -3565 981 -3561
rect 998 -3565 1002 -3561
rect 696 -3735 700 -3731
rect 717 -3735 721 -3731
rect 653 -3766 657 -3762
rect 674 -3766 678 -3762
rect 684 -3984 688 -3980
rect 705 -3984 709 -3980
rect 641 -4015 645 -4011
rect 662 -4015 666 -4011
<< nsubstratencontact >>
rect 1059 1708 1063 1712
rect 1076 1708 1080 1712
rect 903 1681 907 1685
rect 920 1681 924 1685
rect 859 1651 863 1655
rect 859 1634 863 1638
rect 994 1665 998 1669
rect 1011 1665 1015 1669
rect 859 1600 863 1604
rect 1168 1696 1172 1700
rect 1185 1696 1189 1700
rect 1195 1696 1199 1700
rect 1212 1696 1216 1700
rect 3107 1681 3111 1685
rect 3124 1681 3128 1685
rect 2951 1654 2955 1658
rect 2968 1654 2972 1658
rect 859 1583 863 1587
rect 1108 1571 1112 1575
rect 1125 1571 1129 1575
rect 1230 1626 1234 1630
rect 1247 1626 1251 1630
rect 2907 1624 2911 1628
rect 2907 1607 2911 1611
rect 3042 1638 3046 1642
rect 3059 1638 3063 1642
rect 2907 1573 2911 1577
rect 3216 1669 3220 1673
rect 3233 1669 3237 1673
rect 3243 1669 3247 1673
rect 3260 1669 3264 1673
rect 2907 1556 2911 1560
rect 3156 1544 3160 1548
rect 3173 1544 3177 1548
rect 3278 1599 3282 1603
rect 3295 1599 3299 1603
rect -1334 415 -1330 419
rect -1312 415 -1308 419
rect -1302 415 -1298 419
rect -1280 415 -1276 419
rect 3961 412 3965 416
rect 3983 412 3987 416
rect 3993 412 3997 416
rect 4015 412 4019 416
rect -1535 407 -1531 411
rect -1513 407 -1509 411
rect -1483 407 -1479 411
rect -1461 407 -1457 411
rect -1431 407 -1427 411
rect -1409 407 -1405 411
rect -1379 407 -1375 411
rect -1357 407 -1353 411
rect 3760 404 3764 408
rect 3782 404 3786 408
rect 3812 404 3816 408
rect 3834 404 3838 408
rect 3864 404 3868 408
rect 3886 404 3890 408
rect 3916 404 3920 408
rect 3938 404 3942 408
rect 1613 109 1617 113
rect 1635 109 1639 113
rect 1645 109 1649 113
rect 1667 109 1671 113
rect 1412 101 1416 105
rect 1434 101 1438 105
rect 1464 101 1468 105
rect 1486 101 1490 105
rect 1516 101 1520 105
rect 1538 101 1542 105
rect 1568 101 1572 105
rect 1590 101 1594 105
rect 1162 43 1166 47
rect 1179 43 1183 47
rect -208 14 -204 18
rect -186 14 -182 18
rect -176 14 -172 18
rect -154 14 -150 18
rect 1118 13 1122 17
rect -409 6 -405 10
rect -387 6 -383 10
rect -357 6 -353 10
rect -335 6 -331 10
rect -305 6 -301 10
rect -283 6 -279 10
rect -253 6 -249 10
rect -231 6 -227 10
rect 1118 -4 1122 0
rect 1118 -38 1122 -34
rect 811 -53 815 -49
rect 828 -53 832 -49
rect 1118 -55 1122 -51
rect 441 -138 445 -134
rect 458 -138 462 -134
rect 468 -138 472 -134
rect 485 -138 489 -134
rect 249 -156 253 -152
rect 266 -156 270 -152
rect 205 -186 209 -182
rect 205 -203 209 -199
rect 205 -237 209 -233
rect -212 -241 -208 -237
rect -190 -241 -186 -237
rect -180 -241 -176 -237
rect -158 -241 -154 -237
rect -413 -249 -409 -245
rect -391 -249 -387 -245
rect -361 -249 -357 -245
rect -339 -249 -335 -245
rect -309 -249 -305 -245
rect -287 -249 -283 -245
rect -257 -249 -253 -245
rect -235 -249 -231 -245
rect 205 -254 209 -250
rect 503 -208 507 -204
rect 520 -208 524 -204
rect 1628 -167 1632 -163
rect 1650 -167 1654 -163
rect 1660 -167 1664 -163
rect 1682 -167 1686 -163
rect 1157 -177 1161 -173
rect 1174 -177 1178 -173
rect 1427 -175 1431 -171
rect 1449 -175 1453 -171
rect 1479 -175 1483 -171
rect 1501 -175 1505 -171
rect 1531 -175 1535 -171
rect 1553 -175 1557 -171
rect 1583 -175 1587 -171
rect 1605 -175 1609 -171
rect 860 -190 864 -186
rect 877 -190 881 -186
rect 1113 -207 1117 -203
rect 1113 -224 1117 -220
rect 166 -300 170 -296
rect 183 -300 187 -296
rect 193 -300 197 -296
rect 210 -300 214 -296
rect 1113 -258 1117 -254
rect 1113 -275 1117 -271
rect 228 -370 232 -366
rect 245 -370 249 -366
rect 955 -700 959 -696
rect 972 -700 976 -696
rect 1206 -702 1210 -698
rect 1223 -702 1227 -698
rect 621 -789 625 -785
rect 638 -789 642 -785
rect 648 -789 652 -785
rect 665 -789 669 -785
rect -115 -823 -111 -819
rect -93 -823 -89 -819
rect -83 -823 -79 -819
rect -61 -823 -57 -819
rect -316 -831 -312 -827
rect -294 -831 -290 -827
rect -264 -831 -260 -827
rect -242 -831 -238 -827
rect -212 -831 -208 -827
rect -190 -831 -186 -827
rect -160 -831 -156 -827
rect -138 -831 -134 -827
rect 683 -859 687 -855
rect 700 -859 704 -855
rect 1004 -837 1008 -833
rect 1021 -837 1025 -833
rect 237 -942 241 -938
rect 254 -942 258 -938
rect 193 -972 197 -968
rect 193 -989 197 -985
rect 1255 -839 1259 -835
rect 1272 -839 1276 -835
rect 2012 -840 2016 -836
rect 2034 -840 2038 -836
rect 2044 -840 2048 -836
rect 2066 -840 2070 -836
rect 1811 -848 1815 -844
rect 1833 -848 1837 -844
rect 1863 -848 1867 -844
rect 1885 -848 1889 -844
rect 1915 -848 1919 -844
rect 1937 -848 1941 -844
rect 1967 -848 1971 -844
rect 1989 -848 1993 -844
rect 1609 -907 1613 -903
rect 1626 -907 1630 -903
rect 1565 -937 1569 -933
rect 1565 -954 1569 -950
rect 1565 -988 1569 -984
rect 193 -1023 197 -1019
rect 1565 -1005 1569 -1001
rect 544 -1034 548 -1030
rect 561 -1034 565 -1030
rect 571 -1034 575 -1030
rect 588 -1034 592 -1030
rect 762 -1034 766 -1030
rect 779 -1034 783 -1030
rect 789 -1034 793 -1030
rect 806 -1034 810 -1030
rect 193 -1040 197 -1036
rect -134 -1046 -130 -1042
rect -112 -1046 -108 -1042
rect -102 -1046 -98 -1042
rect -80 -1046 -76 -1042
rect -335 -1054 -331 -1050
rect -313 -1054 -309 -1050
rect -283 -1054 -279 -1050
rect -261 -1054 -257 -1050
rect -231 -1054 -227 -1050
rect -209 -1054 -205 -1050
rect -179 -1054 -175 -1050
rect -157 -1054 -153 -1050
rect 154 -1086 158 -1082
rect 171 -1086 175 -1082
rect 181 -1086 185 -1082
rect 198 -1086 202 -1082
rect -3294 -1149 -3290 -1145
rect -3277 -1149 -3273 -1145
rect -3450 -1176 -3446 -1172
rect -3433 -1176 -3429 -1172
rect -3494 -1206 -3490 -1202
rect -3494 -1223 -3490 -1219
rect -3359 -1192 -3355 -1188
rect -3342 -1192 -3338 -1188
rect -3494 -1257 -3490 -1253
rect -3185 -1161 -3181 -1157
rect -3168 -1161 -3164 -1157
rect -3158 -1161 -3154 -1157
rect -3141 -1161 -3137 -1157
rect -3494 -1274 -3490 -1270
rect -3245 -1286 -3241 -1282
rect -3228 -1286 -3224 -1282
rect 216 -1156 220 -1152
rect 233 -1156 237 -1152
rect 606 -1104 610 -1100
rect 623 -1104 627 -1100
rect 824 -1104 828 -1100
rect 841 -1104 845 -1100
rect -3123 -1231 -3119 -1227
rect -3106 -1231 -3102 -1227
rect 556 -1349 560 -1345
rect 573 -1349 577 -1345
rect 583 -1349 587 -1345
rect 600 -1349 604 -1345
rect -134 -1384 -130 -1380
rect -112 -1384 -108 -1380
rect -102 -1384 -98 -1380
rect -80 -1384 -76 -1380
rect -335 -1392 -331 -1388
rect -313 -1392 -309 -1388
rect -283 -1392 -279 -1388
rect -261 -1392 -257 -1388
rect -231 -1392 -227 -1388
rect -209 -1392 -205 -1388
rect -179 -1392 -175 -1388
rect -157 -1392 -153 -1388
rect 618 -1419 622 -1415
rect 635 -1419 639 -1415
rect 1075 -1425 1079 -1421
rect 1092 -1425 1096 -1421
rect 793 -1579 797 -1575
rect 810 -1579 814 -1575
rect 820 -1579 824 -1575
rect 837 -1579 841 -1575
rect 246 -1602 250 -1598
rect 263 -1602 267 -1598
rect 202 -1632 206 -1628
rect 202 -1649 206 -1645
rect 557 -1632 561 -1628
rect 574 -1632 578 -1628
rect 584 -1632 588 -1628
rect 601 -1632 605 -1628
rect 202 -1683 206 -1679
rect 1124 -1562 1128 -1558
rect 1141 -1562 1145 -1558
rect 1372 -1578 1376 -1574
rect 1389 -1578 1393 -1574
rect 202 -1700 206 -1696
rect -149 -1721 -145 -1717
rect -127 -1721 -123 -1717
rect -117 -1721 -113 -1717
rect -95 -1721 -91 -1717
rect -350 -1729 -346 -1725
rect -328 -1729 -324 -1725
rect -298 -1729 -294 -1725
rect -276 -1729 -272 -1725
rect -246 -1729 -242 -1725
rect -224 -1729 -220 -1725
rect -194 -1729 -190 -1725
rect -172 -1729 -168 -1725
rect 163 -1746 167 -1742
rect 180 -1746 184 -1742
rect 190 -1746 194 -1742
rect 207 -1746 211 -1742
rect 619 -1702 623 -1698
rect 636 -1702 640 -1698
rect 855 -1649 859 -1645
rect 872 -1649 876 -1645
rect 2201 -1590 2205 -1586
rect 2223 -1590 2227 -1586
rect 2233 -1590 2237 -1586
rect 2255 -1590 2259 -1586
rect 2000 -1598 2004 -1594
rect 2022 -1598 2026 -1594
rect 2052 -1598 2056 -1594
rect 2074 -1598 2078 -1594
rect 2104 -1598 2108 -1594
rect 2126 -1598 2130 -1594
rect 2156 -1598 2160 -1594
rect 2178 -1598 2182 -1594
rect 1790 -1643 1794 -1639
rect 1807 -1643 1811 -1639
rect 1746 -1673 1750 -1669
rect 1086 -1725 1090 -1721
rect 1103 -1725 1107 -1721
rect 225 -1816 229 -1812
rect 242 -1816 246 -1812
rect 802 -1790 806 -1786
rect 819 -1790 823 -1786
rect 829 -1790 833 -1786
rect 846 -1790 850 -1786
rect 1746 -1690 1750 -1686
rect 1421 -1715 1425 -1711
rect 1438 -1715 1442 -1711
rect 1746 -1724 1750 -1720
rect 1746 -1741 1750 -1737
rect 553 -1903 557 -1899
rect 570 -1903 574 -1899
rect 580 -1903 584 -1899
rect 597 -1903 601 -1899
rect 864 -1860 868 -1856
rect 881 -1860 885 -1856
rect 615 -1973 619 -1969
rect 632 -1973 636 -1969
rect 1135 -1862 1139 -1858
rect 1152 -1862 1156 -1858
rect 541 -2152 545 -2148
rect 558 -2152 562 -2148
rect 568 -2152 572 -2148
rect 585 -2152 589 -2148
rect 603 -2222 607 -2218
rect 620 -2222 624 -2218
rect -149 -2328 -145 -2324
rect -127 -2328 -123 -2324
rect -117 -2328 -113 -2324
rect -95 -2328 -91 -2324
rect -350 -2336 -346 -2332
rect -328 -2336 -324 -2332
rect -298 -2336 -294 -2332
rect -276 -2336 -272 -2332
rect -246 -2336 -242 -2332
rect -224 -2336 -220 -2332
rect -194 -2336 -190 -2332
rect -172 -2336 -168 -2332
rect 243 -2477 247 -2473
rect 260 -2477 264 -2473
rect 199 -2507 203 -2503
rect 199 -2524 203 -2520
rect 1299 -2492 1303 -2488
rect 1316 -2492 1320 -2488
rect 634 -2499 638 -2495
rect 651 -2499 655 -2495
rect 661 -2499 665 -2495
rect 678 -2499 682 -2495
rect 199 -2558 203 -2554
rect 199 -2575 203 -2571
rect 969 -2551 973 -2547
rect 986 -2551 990 -2547
rect 996 -2551 1000 -2547
rect 1013 -2551 1017 -2547
rect -149 -2598 -145 -2594
rect -127 -2598 -123 -2594
rect -117 -2598 -113 -2594
rect -95 -2598 -91 -2594
rect -350 -2606 -346 -2602
rect -328 -2606 -324 -2602
rect -298 -2606 -294 -2602
rect -276 -2606 -272 -2602
rect -246 -2606 -242 -2602
rect -224 -2606 -220 -2602
rect -194 -2606 -190 -2602
rect -172 -2606 -168 -2602
rect 160 -2621 164 -2617
rect 177 -2621 181 -2617
rect 187 -2621 191 -2617
rect 204 -2621 208 -2617
rect 696 -2569 700 -2565
rect 713 -2569 717 -2565
rect 222 -2691 226 -2687
rect 239 -2691 243 -2687
rect 1031 -2621 1035 -2617
rect 1048 -2621 1052 -2617
rect 1348 -2629 1352 -2625
rect 1365 -2629 1369 -2625
rect 635 -2782 639 -2778
rect 652 -2782 656 -2778
rect 662 -2782 666 -2778
rect 679 -2782 683 -2778
rect 1803 -2806 1807 -2802
rect 1820 -2806 1824 -2802
rect 970 -2834 974 -2830
rect 987 -2834 991 -2830
rect 997 -2834 1001 -2830
rect 1014 -2834 1018 -2830
rect 697 -2852 701 -2848
rect 714 -2852 718 -2848
rect 1306 -2881 1310 -2877
rect 1323 -2881 1327 -2877
rect 1032 -2904 1036 -2900
rect 1049 -2904 1053 -2900
rect 2275 -2832 2279 -2828
rect 2297 -2832 2301 -2828
rect 2307 -2832 2311 -2828
rect 2329 -2832 2333 -2828
rect 2074 -2840 2078 -2836
rect 2096 -2840 2100 -2836
rect 2126 -2840 2130 -2836
rect 2148 -2840 2152 -2836
rect 2178 -2840 2182 -2836
rect 2200 -2840 2204 -2836
rect 2230 -2840 2234 -2836
rect 2252 -2840 2256 -2836
rect 631 -3053 635 -3049
rect 648 -3053 652 -3049
rect 658 -3053 662 -3049
rect 675 -3053 679 -3049
rect 1355 -3018 1359 -3014
rect 1372 -3018 1376 -3014
rect 1852 -2943 1856 -2939
rect 1869 -2943 1873 -2939
rect 1598 -3037 1602 -3033
rect 1615 -3037 1619 -3033
rect 693 -3123 697 -3119
rect 710 -3123 714 -3119
rect 1300 -3236 1304 -3232
rect 1317 -3236 1321 -3232
rect 1327 -3236 1331 -3232
rect 1344 -3236 1348 -3232
rect 1647 -3174 1651 -3170
rect 1664 -3174 1668 -3170
rect 619 -3302 623 -3298
rect 636 -3302 640 -3298
rect 646 -3302 650 -3298
rect 663 -3302 667 -3298
rect 960 -3368 964 -3364
rect 977 -3368 981 -3364
rect 987 -3368 991 -3364
rect 1004 -3368 1008 -3364
rect 681 -3372 685 -3368
rect 698 -3372 702 -3368
rect 1362 -3306 1366 -3302
rect 1379 -3306 1383 -3302
rect 1022 -3438 1026 -3434
rect 1039 -3438 1043 -3434
rect 636 -3569 640 -3565
rect 653 -3569 657 -3565
rect 663 -3569 667 -3565
rect 680 -3569 684 -3565
rect 698 -3639 702 -3635
rect 715 -3639 719 -3635
rect 624 -3818 628 -3814
rect 641 -3818 645 -3814
rect 651 -3818 655 -3814
rect 668 -3818 672 -3814
rect 686 -3888 690 -3884
rect 703 -3888 707 -3884
<< polysilicon >>
rect 1069 1701 1071 1704
rect 797 1673 879 1675
rect 913 1674 915 1677
rect 877 1651 879 1673
rect 771 1643 774 1645
rect 794 1643 812 1645
rect 852 1643 855 1645
rect 1004 1658 1006 1661
rect 877 1628 879 1631
rect 797 1621 879 1623
rect 877 1618 879 1621
rect 913 1616 915 1634
rect 1178 1689 1180 1692
rect 1205 1689 1207 1692
rect 3117 1674 3119 1677
rect 877 1595 879 1598
rect 1004 1600 1006 1618
rect 1069 1615 1071 1621
rect 1178 1621 1180 1649
rect 1205 1637 1207 1649
rect 2845 1646 2927 1648
rect 2961 1647 2963 1650
rect 1205 1635 1215 1637
rect 1178 1619 1199 1621
rect 1197 1615 1199 1619
rect 1069 1613 1089 1615
rect 1069 1601 1071 1604
rect 771 1592 774 1594
rect 794 1592 812 1594
rect 852 1592 855 1594
rect 913 1593 915 1596
rect 1004 1577 1006 1580
rect 1069 1515 1071 1521
rect 1054 1513 1071 1515
rect 1054 1496 1056 1513
rect 1087 1496 1089 1613
rect 1197 1571 1199 1575
rect 1118 1564 1120 1567
rect 1213 1558 1215 1635
rect 2925 1624 2927 1646
rect 1240 1619 1242 1622
rect 2819 1616 2822 1618
rect 2842 1616 2860 1618
rect 2900 1616 2903 1618
rect 3052 1631 3054 1634
rect 2925 1601 2927 1604
rect 2845 1594 2927 1596
rect 2925 1591 2927 1594
rect 1240 1561 1242 1579
rect 2961 1589 2963 1607
rect 3226 1662 3228 1665
rect 3253 1662 3255 1665
rect 2925 1568 2927 1571
rect 3052 1573 3054 1591
rect 3117 1588 3119 1594
rect 3226 1594 3228 1622
rect 3253 1610 3255 1622
rect 3253 1608 3263 1610
rect 3226 1592 3247 1594
rect 3245 1588 3247 1592
rect 3117 1586 3137 1588
rect 3117 1574 3119 1577
rect 2819 1565 2822 1567
rect 2842 1565 2860 1567
rect 2900 1565 2903 1567
rect 2961 1566 2963 1569
rect 1197 1556 1215 1558
rect 1197 1550 1199 1556
rect 1118 1506 1120 1524
rect 3052 1550 3054 1553
rect 1240 1538 1242 1541
rect 1197 1507 1199 1510
rect 3117 1488 3119 1494
rect 1118 1483 1120 1486
rect 3102 1486 3119 1488
rect 1054 1473 1056 1476
rect 1087 1473 1089 1476
rect 3102 1469 3104 1486
rect 3135 1469 3137 1586
rect 3245 1544 3247 1548
rect 3166 1537 3168 1540
rect 3261 1531 3263 1608
rect 3288 1592 3290 1595
rect 3288 1534 3290 1552
rect 3245 1529 3263 1531
rect 3245 1523 3247 1529
rect 3166 1479 3168 1497
rect 3288 1511 3290 1514
rect 3245 1480 3247 1483
rect 3166 1456 3168 1459
rect 3102 1446 3104 1449
rect 3135 1446 3137 1449
rect -1322 407 -1320 411
rect -1290 407 -1288 411
rect -1523 399 -1521 403
rect -1471 399 -1469 403
rect -1419 399 -1417 403
rect -1367 399 -1365 403
rect 3973 404 3975 408
rect 4005 404 4007 408
rect 3772 396 3774 400
rect 3824 396 3826 400
rect 3876 396 3878 400
rect 3928 396 3930 400
rect -1523 350 -1521 359
rect -1471 350 -1469 359
rect -1419 350 -1417 359
rect -1367 350 -1365 359
rect -1322 347 -1320 367
rect -1290 347 -1288 367
rect 3772 347 3774 356
rect 3824 347 3826 356
rect 3876 347 3878 356
rect 3928 347 3930 356
rect -1523 337 -1521 341
rect -1471 337 -1469 341
rect -1419 323 -1417 332
rect -1367 323 -1365 332
rect 3973 344 3975 364
rect 4005 344 4007 364
rect 3772 334 3774 338
rect 3824 334 3826 338
rect -1322 323 -1320 327
rect -1290 323 -1288 327
rect -1419 300 -1417 303
rect -1367 300 -1365 303
rect -1523 288 -1521 297
rect -1471 288 -1469 297
rect 3876 320 3878 329
rect 3928 320 3930 329
rect 3973 320 3975 324
rect 4005 320 4007 324
rect 3876 297 3878 300
rect 3928 297 3930 300
rect 3772 285 3774 294
rect 3824 285 3826 294
rect -1523 276 -1521 284
rect -1471 276 -1469 284
rect -1419 276 -1417 284
rect -1367 276 -1365 284
rect 3772 273 3774 281
rect 3824 273 3826 281
rect 3876 273 3878 281
rect 3928 273 3930 281
rect -1523 252 -1521 256
rect -1471 252 -1469 256
rect -1419 252 -1417 256
rect -1367 252 -1365 256
rect 3772 249 3774 253
rect 3824 249 3826 253
rect 3876 249 3878 253
rect 3928 249 3930 253
rect 1625 101 1627 105
rect 1657 101 1659 105
rect 1424 93 1426 97
rect 1476 93 1478 97
rect 1528 93 1530 97
rect 1580 93 1582 97
rect 1424 44 1426 53
rect 1476 44 1478 53
rect 1528 44 1530 53
rect 1580 44 1582 53
rect 1625 41 1627 61
rect 1657 41 1659 61
rect 1056 35 1138 37
rect 1172 36 1174 39
rect 1136 13 1138 35
rect -196 6 -194 10
rect -164 6 -162 10
rect -397 -2 -395 2
rect -345 -2 -343 2
rect -293 -2 -291 2
rect -241 -2 -239 2
rect 1030 5 1033 7
rect 1053 5 1071 7
rect 1111 5 1114 7
rect 1424 31 1426 35
rect 1476 31 1478 35
rect 1136 -10 1138 -7
rect 1056 -17 1138 -15
rect 1136 -20 1138 -17
rect -397 -51 -395 -42
rect -345 -51 -343 -42
rect -293 -51 -291 -42
rect -241 -51 -239 -42
rect -196 -54 -194 -34
rect -164 -54 -162 -34
rect 1172 -22 1174 -4
rect 1528 17 1530 26
rect 1580 17 1582 26
rect 1625 17 1627 21
rect 1657 17 1659 21
rect 1528 -6 1530 -3
rect 1580 -6 1582 -3
rect 1424 -18 1426 -9
rect 1476 -18 1478 -9
rect 1136 -43 1138 -40
rect 1424 -30 1426 -22
rect 1476 -30 1478 -22
rect 1528 -30 1530 -22
rect 1580 -30 1582 -22
rect 1030 -46 1033 -44
rect 1053 -46 1071 -44
rect 1111 -46 1114 -44
rect 1172 -45 1174 -42
rect -397 -64 -395 -60
rect -345 -64 -343 -60
rect -293 -78 -291 -69
rect -241 -78 -239 -69
rect 1424 -54 1426 -50
rect 1476 -54 1478 -50
rect 1528 -54 1530 -50
rect 1580 -54 1582 -50
rect 821 -60 823 -57
rect -196 -78 -194 -74
rect -164 -78 -162 -74
rect -293 -101 -291 -98
rect -241 -101 -239 -98
rect -397 -113 -395 -104
rect -345 -113 -343 -104
rect -397 -125 -395 -117
rect -345 -125 -343 -117
rect -293 -125 -291 -117
rect -241 -125 -239 -117
rect 451 -145 453 -142
rect 478 -145 480 -142
rect -397 -149 -395 -145
rect -345 -149 -343 -145
rect -293 -149 -291 -145
rect -241 -149 -239 -145
rect 143 -164 225 -162
rect 259 -163 261 -160
rect 223 -186 225 -164
rect 117 -194 120 -192
rect 140 -194 158 -192
rect 198 -194 201 -192
rect 821 -146 823 -140
rect 821 -148 841 -146
rect 821 -160 823 -157
rect 223 -209 225 -206
rect 143 -216 225 -214
rect 223 -219 225 -216
rect 259 -221 261 -203
rect 451 -213 453 -185
rect 478 -197 480 -185
rect 478 -199 488 -197
rect 451 -215 472 -213
rect 470 -219 472 -215
rect 223 -242 225 -239
rect 117 -245 120 -243
rect 140 -245 158 -243
rect 198 -245 201 -243
rect 259 -244 261 -241
rect -200 -249 -198 -245
rect -168 -249 -166 -245
rect -401 -257 -399 -253
rect -349 -257 -347 -253
rect -297 -257 -295 -253
rect -245 -257 -243 -253
rect 470 -263 472 -259
rect 486 -276 488 -199
rect 513 -215 515 -212
rect 821 -246 823 -240
rect 806 -248 823 -246
rect 513 -273 515 -255
rect 806 -265 808 -248
rect 839 -265 841 -148
rect 1640 -175 1642 -171
rect 1672 -175 1674 -171
rect 1051 -185 1133 -183
rect 1167 -184 1169 -181
rect 1439 -183 1441 -179
rect 1491 -183 1493 -179
rect 1543 -183 1545 -179
rect 1595 -183 1597 -179
rect 870 -197 872 -194
rect 1131 -207 1133 -185
rect 1025 -215 1028 -213
rect 1048 -215 1066 -213
rect 1106 -215 1109 -213
rect 1131 -230 1133 -227
rect 1051 -237 1133 -235
rect 870 -255 872 -237
rect 1131 -240 1133 -237
rect 470 -278 488 -276
rect 470 -284 472 -278
rect -401 -306 -399 -297
rect -349 -306 -347 -297
rect -297 -306 -295 -297
rect -245 -306 -243 -297
rect -200 -309 -198 -289
rect -168 -309 -166 -289
rect 176 -307 178 -304
rect 203 -307 205 -304
rect -401 -319 -399 -315
rect -349 -319 -347 -315
rect -297 -333 -295 -324
rect -245 -333 -243 -324
rect -200 -333 -198 -329
rect -168 -333 -166 -329
rect 1167 -242 1169 -224
rect 1439 -232 1441 -223
rect 1491 -232 1493 -223
rect 1543 -232 1545 -223
rect 1595 -232 1597 -223
rect 1640 -235 1642 -215
rect 1672 -235 1674 -215
rect 1131 -263 1133 -260
rect 1439 -245 1441 -241
rect 1491 -245 1493 -241
rect 1025 -266 1028 -264
rect 1048 -266 1066 -264
rect 1106 -266 1109 -264
rect 1167 -265 1169 -262
rect 870 -278 872 -275
rect 806 -288 808 -285
rect 839 -288 841 -285
rect 1543 -259 1545 -250
rect 1595 -259 1597 -250
rect 1640 -259 1642 -255
rect 1672 -259 1674 -255
rect 1543 -282 1545 -279
rect 1595 -282 1597 -279
rect 513 -296 515 -293
rect 1439 -294 1441 -285
rect 1491 -294 1493 -285
rect 1439 -306 1441 -298
rect 1491 -306 1493 -298
rect 1543 -306 1545 -298
rect 1595 -306 1597 -298
rect 470 -327 472 -324
rect 1439 -330 1441 -326
rect 1491 -330 1493 -326
rect 1543 -330 1545 -326
rect 1595 -330 1597 -326
rect -297 -356 -295 -353
rect -245 -356 -243 -353
rect -401 -368 -399 -359
rect -349 -368 -347 -359
rect -401 -380 -399 -372
rect -349 -380 -347 -372
rect -297 -380 -295 -372
rect -245 -380 -243 -372
rect 176 -375 178 -347
rect 203 -359 205 -347
rect 203 -361 213 -359
rect 176 -377 197 -375
rect 195 -381 197 -377
rect -401 -404 -399 -400
rect -349 -404 -347 -400
rect -297 -404 -295 -400
rect -245 -404 -243 -400
rect 195 -425 197 -421
rect 211 -438 213 -361
rect 238 -377 240 -374
rect 238 -435 240 -417
rect 195 -440 213 -438
rect 195 -446 197 -440
rect 238 -458 240 -455
rect 195 -489 197 -486
rect 965 -707 967 -704
rect 1216 -709 1218 -706
rect 631 -796 633 -793
rect 658 -796 660 -793
rect 965 -793 967 -787
rect 965 -795 985 -793
rect -103 -831 -101 -827
rect -71 -831 -69 -827
rect -304 -839 -302 -835
rect -252 -839 -250 -835
rect -200 -839 -198 -835
rect -148 -839 -146 -835
rect 965 -807 967 -804
rect 631 -864 633 -836
rect 658 -848 660 -836
rect 658 -850 668 -848
rect 631 -866 652 -864
rect 650 -870 652 -866
rect -304 -888 -302 -879
rect -252 -888 -250 -879
rect -200 -888 -198 -879
rect -148 -888 -146 -879
rect -103 -891 -101 -871
rect -71 -891 -69 -871
rect -304 -901 -302 -897
rect -252 -901 -250 -897
rect -200 -915 -198 -906
rect -148 -915 -146 -906
rect -103 -915 -101 -911
rect -71 -915 -69 -911
rect 650 -914 652 -910
rect 666 -927 668 -850
rect 693 -866 695 -863
rect 965 -893 967 -887
rect 950 -895 967 -893
rect 693 -924 695 -906
rect 950 -912 952 -895
rect 983 -912 985 -795
rect 1216 -795 1218 -789
rect 1216 -797 1236 -795
rect 1216 -809 1218 -806
rect 1014 -844 1016 -841
rect 1014 -902 1016 -884
rect 1216 -895 1218 -889
rect 1201 -897 1218 -895
rect 650 -929 668 -927
rect 650 -935 652 -929
rect -200 -938 -198 -935
rect -148 -938 -146 -935
rect -304 -950 -302 -941
rect -252 -950 -250 -941
rect 131 -950 213 -948
rect 247 -949 249 -946
rect -304 -962 -302 -954
rect -252 -962 -250 -954
rect -200 -962 -198 -954
rect -148 -962 -146 -954
rect 211 -972 213 -950
rect 105 -980 108 -978
rect 128 -980 146 -978
rect 186 -980 189 -978
rect -304 -986 -302 -982
rect -252 -986 -250 -982
rect -200 -986 -198 -982
rect -148 -986 -146 -982
rect 1201 -914 1203 -897
rect 1234 -914 1236 -797
rect 1265 -846 1267 -843
rect 2024 -848 2026 -844
rect 2056 -848 2058 -844
rect 1823 -856 1825 -852
rect 1875 -856 1877 -852
rect 1927 -856 1929 -852
rect 1979 -856 1981 -852
rect 1265 -904 1267 -886
rect 1014 -925 1016 -922
rect 950 -935 952 -932
rect 983 -935 985 -932
rect 1823 -905 1825 -896
rect 1875 -905 1877 -896
rect 1927 -905 1929 -896
rect 1979 -905 1981 -896
rect 2024 -908 2026 -888
rect 2056 -908 2058 -888
rect 1503 -915 1585 -913
rect 1619 -914 1621 -911
rect 1265 -927 1267 -924
rect 1201 -937 1203 -934
rect 1234 -937 1236 -934
rect 1583 -937 1585 -915
rect 693 -947 695 -944
rect 1477 -945 1480 -943
rect 1500 -945 1518 -943
rect 1558 -945 1561 -943
rect 1823 -918 1825 -914
rect 1875 -918 1877 -914
rect 1583 -960 1585 -957
rect 1503 -967 1585 -965
rect 1583 -970 1585 -967
rect 650 -978 652 -975
rect 211 -995 213 -992
rect 131 -1002 213 -1000
rect 211 -1005 213 -1002
rect 247 -1007 249 -989
rect 1619 -972 1621 -954
rect 1927 -932 1929 -923
rect 1979 -932 1981 -923
rect 2024 -932 2026 -928
rect 2056 -932 2058 -928
rect 1927 -955 1929 -952
rect 1979 -955 1981 -952
rect 1823 -967 1825 -958
rect 1875 -967 1877 -958
rect 1583 -993 1585 -990
rect 1823 -979 1825 -971
rect 1875 -979 1877 -971
rect 1927 -979 1929 -971
rect 1979 -979 1981 -971
rect 1477 -996 1480 -994
rect 1500 -996 1518 -994
rect 1558 -996 1561 -994
rect 1619 -995 1621 -992
rect 1823 -1003 1825 -999
rect 1875 -1003 1877 -999
rect 1927 -1003 1929 -999
rect 1979 -1003 1981 -999
rect 211 -1028 213 -1025
rect 105 -1031 108 -1029
rect 128 -1031 146 -1029
rect 186 -1031 189 -1029
rect 247 -1030 249 -1027
rect 554 -1041 556 -1038
rect 581 -1041 583 -1038
rect 772 -1041 774 -1038
rect 799 -1041 801 -1038
rect -122 -1054 -120 -1050
rect -90 -1054 -88 -1050
rect -323 -1062 -321 -1058
rect -271 -1062 -269 -1058
rect -219 -1062 -217 -1058
rect -167 -1062 -165 -1058
rect 164 -1093 166 -1090
rect 191 -1093 193 -1090
rect -323 -1111 -321 -1102
rect -271 -1111 -269 -1102
rect -219 -1111 -217 -1102
rect -167 -1111 -165 -1102
rect -122 -1114 -120 -1094
rect -90 -1114 -88 -1094
rect -323 -1124 -321 -1120
rect -271 -1124 -269 -1120
rect -3284 -1156 -3282 -1153
rect -3556 -1184 -3474 -1182
rect -3440 -1183 -3438 -1180
rect -3476 -1206 -3474 -1184
rect -3582 -1214 -3579 -1212
rect -3559 -1214 -3541 -1212
rect -3501 -1214 -3498 -1212
rect -3349 -1199 -3347 -1196
rect -3476 -1229 -3474 -1226
rect -3556 -1236 -3474 -1234
rect -3476 -1239 -3474 -1236
rect -3440 -1241 -3438 -1223
rect -219 -1138 -217 -1129
rect -167 -1138 -165 -1129
rect 554 -1109 556 -1081
rect 581 -1093 583 -1081
rect 581 -1095 591 -1093
rect 554 -1111 575 -1109
rect 573 -1115 575 -1111
rect -122 -1138 -120 -1134
rect -90 -1138 -88 -1134
rect -219 -1161 -217 -1158
rect -167 -1161 -165 -1158
rect 164 -1161 166 -1133
rect 191 -1145 193 -1133
rect 191 -1147 201 -1145
rect 164 -1163 185 -1161
rect -3175 -1168 -3173 -1165
rect -3148 -1168 -3146 -1165
rect -323 -1173 -321 -1164
rect -271 -1173 -269 -1164
rect 183 -1167 185 -1163
rect -323 -1185 -321 -1177
rect -271 -1185 -269 -1177
rect -219 -1185 -217 -1177
rect -167 -1185 -165 -1177
rect -3476 -1262 -3474 -1259
rect -3349 -1257 -3347 -1239
rect -3284 -1242 -3282 -1236
rect -3175 -1236 -3173 -1208
rect -3148 -1220 -3146 -1208
rect -323 -1209 -321 -1205
rect -271 -1209 -269 -1205
rect -219 -1209 -217 -1205
rect -167 -1209 -165 -1205
rect 183 -1211 185 -1207
rect -3148 -1222 -3138 -1220
rect -3175 -1238 -3154 -1236
rect -3156 -1242 -3154 -1238
rect -3284 -1244 -3264 -1242
rect -3284 -1256 -3282 -1253
rect -3582 -1265 -3579 -1263
rect -3559 -1265 -3541 -1263
rect -3501 -1265 -3498 -1263
rect -3440 -1264 -3438 -1261
rect -3349 -1280 -3347 -1277
rect -3284 -1342 -3282 -1336
rect -3299 -1344 -3282 -1342
rect -3299 -1361 -3297 -1344
rect -3266 -1361 -3264 -1244
rect -3156 -1286 -3154 -1282
rect -3235 -1293 -3233 -1290
rect -3140 -1299 -3138 -1222
rect 199 -1224 201 -1147
rect 573 -1159 575 -1155
rect 226 -1163 228 -1160
rect 589 -1172 591 -1095
rect 616 -1111 618 -1108
rect 772 -1109 774 -1081
rect 799 -1093 801 -1081
rect 799 -1095 809 -1093
rect 772 -1111 793 -1109
rect 791 -1115 793 -1111
rect 616 -1169 618 -1151
rect 791 -1159 793 -1155
rect 573 -1174 591 -1172
rect 573 -1180 575 -1174
rect 226 -1221 228 -1203
rect 807 -1172 809 -1095
rect 834 -1111 836 -1108
rect 834 -1169 836 -1151
rect 791 -1174 809 -1172
rect 791 -1180 793 -1174
rect 616 -1192 618 -1189
rect 834 -1192 836 -1189
rect 183 -1226 201 -1224
rect 183 -1232 185 -1226
rect -3113 -1238 -3111 -1235
rect 573 -1223 575 -1220
rect 791 -1223 793 -1220
rect 226 -1244 228 -1241
rect 183 -1275 185 -1272
rect -3113 -1296 -3111 -1278
rect -3156 -1301 -3138 -1299
rect -3156 -1307 -3154 -1301
rect -3235 -1351 -3233 -1333
rect -3113 -1319 -3111 -1316
rect -3156 -1350 -3154 -1347
rect 566 -1356 568 -1353
rect 593 -1356 595 -1353
rect -3235 -1374 -3233 -1371
rect -3299 -1384 -3297 -1381
rect -3266 -1384 -3264 -1381
rect -122 -1392 -120 -1388
rect -90 -1392 -88 -1388
rect -323 -1400 -321 -1396
rect -271 -1400 -269 -1396
rect -219 -1400 -217 -1396
rect -167 -1400 -165 -1396
rect 566 -1424 568 -1396
rect 593 -1408 595 -1396
rect 593 -1410 603 -1408
rect 566 -1426 587 -1424
rect 585 -1430 587 -1426
rect -323 -1449 -321 -1440
rect -271 -1449 -269 -1440
rect -219 -1449 -217 -1440
rect -167 -1449 -165 -1440
rect -122 -1452 -120 -1432
rect -90 -1452 -88 -1432
rect -323 -1462 -321 -1458
rect -271 -1462 -269 -1458
rect -219 -1476 -217 -1467
rect -167 -1476 -165 -1467
rect -122 -1476 -120 -1472
rect -90 -1476 -88 -1472
rect 585 -1474 587 -1470
rect 601 -1487 603 -1410
rect 628 -1426 630 -1423
rect 1085 -1432 1087 -1429
rect 628 -1484 630 -1466
rect 585 -1489 603 -1487
rect 585 -1495 587 -1489
rect -219 -1499 -217 -1496
rect -167 -1499 -165 -1496
rect -323 -1511 -321 -1502
rect -271 -1511 -269 -1502
rect -323 -1523 -321 -1515
rect -271 -1523 -269 -1515
rect -219 -1523 -217 -1515
rect -167 -1523 -165 -1515
rect 628 -1507 630 -1504
rect 1085 -1518 1087 -1512
rect 1085 -1520 1105 -1518
rect 1085 -1532 1087 -1529
rect 585 -1538 587 -1535
rect -323 -1547 -321 -1543
rect -271 -1547 -269 -1543
rect -219 -1547 -217 -1543
rect -167 -1547 -165 -1543
rect 803 -1586 805 -1583
rect 830 -1586 832 -1583
rect 140 -1610 222 -1608
rect 256 -1609 258 -1606
rect 220 -1632 222 -1610
rect 114 -1640 117 -1638
rect 137 -1640 155 -1638
rect 195 -1640 198 -1638
rect 1085 -1618 1087 -1612
rect 1070 -1620 1087 -1618
rect 567 -1639 569 -1636
rect 594 -1639 596 -1636
rect 220 -1655 222 -1652
rect 140 -1662 222 -1660
rect 220 -1665 222 -1662
rect 256 -1667 258 -1649
rect 220 -1688 222 -1685
rect 803 -1654 805 -1626
rect 830 -1638 832 -1626
rect 1070 -1637 1072 -1620
rect 1103 -1637 1105 -1520
rect 1134 -1569 1136 -1566
rect 1382 -1585 1384 -1582
rect 1134 -1627 1136 -1609
rect 830 -1640 840 -1638
rect 803 -1656 824 -1654
rect 822 -1660 824 -1656
rect 114 -1691 117 -1689
rect 137 -1691 155 -1689
rect 195 -1691 198 -1689
rect 256 -1690 258 -1687
rect 567 -1707 569 -1679
rect 594 -1691 596 -1679
rect 594 -1693 604 -1691
rect 567 -1709 588 -1707
rect 586 -1713 588 -1709
rect -137 -1729 -135 -1725
rect -105 -1729 -103 -1725
rect -338 -1737 -336 -1733
rect -286 -1737 -284 -1733
rect -234 -1737 -232 -1733
rect -182 -1737 -180 -1733
rect 173 -1753 175 -1750
rect 200 -1753 202 -1750
rect -338 -1786 -336 -1777
rect -286 -1786 -284 -1777
rect -234 -1786 -232 -1777
rect -182 -1786 -180 -1777
rect -137 -1789 -135 -1769
rect -105 -1789 -103 -1769
rect -338 -1799 -336 -1795
rect -286 -1799 -284 -1795
rect -234 -1813 -232 -1804
rect -182 -1813 -180 -1804
rect 586 -1757 588 -1753
rect 602 -1770 604 -1693
rect 822 -1704 824 -1700
rect 629 -1709 631 -1706
rect 838 -1717 840 -1640
rect 865 -1656 867 -1653
rect 1134 -1650 1136 -1647
rect 1070 -1660 1072 -1657
rect 1103 -1660 1105 -1657
rect 2213 -1598 2215 -1594
rect 2245 -1598 2247 -1594
rect 2012 -1606 2014 -1602
rect 2064 -1606 2066 -1602
rect 2116 -1606 2118 -1602
rect 2168 -1606 2170 -1602
rect 1684 -1651 1766 -1649
rect 1800 -1650 1802 -1647
rect 1382 -1671 1384 -1665
rect 1382 -1673 1402 -1671
rect 1764 -1673 1766 -1651
rect 1382 -1685 1384 -1682
rect 865 -1714 867 -1696
rect 822 -1719 840 -1717
rect 822 -1725 824 -1719
rect 629 -1767 631 -1749
rect 1096 -1732 1098 -1729
rect 865 -1737 867 -1734
rect 586 -1772 604 -1770
rect 586 -1778 588 -1772
rect -137 -1813 -135 -1809
rect -105 -1813 -103 -1809
rect 173 -1821 175 -1793
rect 200 -1805 202 -1793
rect 200 -1807 210 -1805
rect 173 -1823 194 -1821
rect 192 -1827 194 -1823
rect -234 -1836 -232 -1833
rect -182 -1836 -180 -1833
rect -338 -1848 -336 -1839
rect -286 -1848 -284 -1839
rect -338 -1860 -336 -1852
rect -286 -1860 -284 -1852
rect -234 -1860 -232 -1852
rect -182 -1860 -180 -1852
rect 192 -1871 194 -1867
rect -338 -1884 -336 -1880
rect -286 -1884 -284 -1880
rect -234 -1884 -232 -1880
rect -182 -1884 -180 -1880
rect 208 -1884 210 -1807
rect 822 -1768 824 -1765
rect 629 -1790 631 -1787
rect 812 -1797 814 -1794
rect 839 -1797 841 -1794
rect 235 -1823 237 -1820
rect 586 -1821 588 -1818
rect 1382 -1771 1384 -1765
rect 1367 -1773 1384 -1771
rect 1367 -1790 1369 -1773
rect 1400 -1790 1402 -1673
rect 1658 -1681 1661 -1679
rect 1681 -1681 1699 -1679
rect 1739 -1681 1742 -1679
rect 2012 -1655 2014 -1646
rect 2064 -1655 2066 -1646
rect 2116 -1655 2118 -1646
rect 2168 -1655 2170 -1646
rect 2213 -1658 2215 -1638
rect 2245 -1658 2247 -1638
rect 2012 -1668 2014 -1664
rect 2064 -1668 2066 -1664
rect 1764 -1696 1766 -1693
rect 1684 -1703 1766 -1701
rect 1764 -1706 1766 -1703
rect 1431 -1722 1433 -1719
rect 1800 -1708 1802 -1690
rect 2116 -1682 2118 -1673
rect 2168 -1682 2170 -1673
rect 2213 -1682 2215 -1678
rect 2245 -1682 2247 -1678
rect 2116 -1705 2118 -1702
rect 2168 -1705 2170 -1702
rect 1764 -1729 1766 -1726
rect 2012 -1717 2014 -1708
rect 2064 -1717 2066 -1708
rect 1658 -1732 1661 -1730
rect 1681 -1732 1699 -1730
rect 1739 -1732 1742 -1730
rect 1800 -1731 1802 -1728
rect 2012 -1729 2014 -1721
rect 2064 -1729 2066 -1721
rect 2116 -1729 2118 -1721
rect 2168 -1729 2170 -1721
rect 2012 -1753 2014 -1749
rect 2064 -1753 2066 -1749
rect 2116 -1753 2118 -1749
rect 2168 -1753 2170 -1749
rect 1431 -1780 1433 -1762
rect 1431 -1803 1433 -1800
rect 1096 -1818 1098 -1812
rect 1367 -1813 1369 -1810
rect 1400 -1813 1402 -1810
rect 1096 -1820 1116 -1818
rect 1096 -1832 1098 -1829
rect 235 -1881 237 -1863
rect 812 -1865 814 -1837
rect 839 -1849 841 -1837
rect 839 -1851 849 -1849
rect 812 -1867 833 -1865
rect 831 -1871 833 -1867
rect 192 -1886 210 -1884
rect 192 -1892 194 -1886
rect 235 -1904 237 -1901
rect 563 -1910 565 -1907
rect 590 -1910 592 -1907
rect 192 -1935 194 -1932
rect 831 -1915 833 -1911
rect 847 -1928 849 -1851
rect 874 -1867 876 -1864
rect 874 -1925 876 -1907
rect 1096 -1918 1098 -1912
rect 1081 -1920 1098 -1918
rect 831 -1930 849 -1928
rect 831 -1936 833 -1930
rect 563 -1978 565 -1950
rect 590 -1962 592 -1950
rect 590 -1964 600 -1962
rect 563 -1980 584 -1978
rect 582 -1984 584 -1980
rect 582 -2028 584 -2024
rect 598 -2041 600 -1964
rect 1081 -1937 1083 -1920
rect 1114 -1937 1116 -1820
rect 1145 -1869 1147 -1866
rect 1145 -1927 1147 -1909
rect 874 -1948 876 -1945
rect 1145 -1950 1147 -1947
rect 1081 -1960 1083 -1957
rect 1114 -1960 1116 -1957
rect 625 -1980 627 -1977
rect 831 -1979 833 -1976
rect 625 -2038 627 -2020
rect 582 -2043 600 -2041
rect 582 -2049 584 -2043
rect 625 -2061 627 -2058
rect 582 -2092 584 -2089
rect 551 -2159 553 -2156
rect 578 -2159 580 -2156
rect 551 -2227 553 -2199
rect 578 -2211 580 -2199
rect 578 -2213 588 -2211
rect 551 -2229 572 -2227
rect 570 -2233 572 -2229
rect 570 -2277 572 -2273
rect 586 -2290 588 -2213
rect 613 -2229 615 -2226
rect 613 -2287 615 -2269
rect 570 -2292 588 -2290
rect 570 -2298 572 -2292
rect -137 -2336 -135 -2332
rect -105 -2336 -103 -2332
rect -338 -2344 -336 -2340
rect -286 -2344 -284 -2340
rect -234 -2344 -232 -2340
rect -182 -2344 -180 -2340
rect 613 -2310 615 -2307
rect 570 -2341 572 -2338
rect -338 -2393 -336 -2384
rect -286 -2393 -284 -2384
rect -234 -2393 -232 -2384
rect -182 -2393 -180 -2384
rect -137 -2396 -135 -2376
rect -105 -2396 -103 -2376
rect -338 -2406 -336 -2402
rect -286 -2406 -284 -2402
rect -234 -2420 -232 -2411
rect -182 -2420 -180 -2411
rect -137 -2420 -135 -2416
rect -105 -2420 -103 -2416
rect -234 -2443 -232 -2440
rect -182 -2443 -180 -2440
rect -338 -2455 -336 -2446
rect -286 -2455 -284 -2446
rect -338 -2467 -336 -2459
rect -286 -2467 -284 -2459
rect -234 -2467 -232 -2459
rect -182 -2467 -180 -2459
rect 137 -2485 219 -2483
rect 253 -2484 255 -2481
rect -338 -2491 -336 -2487
rect -286 -2491 -284 -2487
rect -234 -2491 -232 -2487
rect -182 -2491 -180 -2487
rect 217 -2507 219 -2485
rect 111 -2515 114 -2513
rect 134 -2515 152 -2513
rect 192 -2515 195 -2513
rect 1309 -2499 1311 -2496
rect 644 -2506 646 -2503
rect 671 -2506 673 -2503
rect 217 -2530 219 -2527
rect 137 -2537 219 -2535
rect 217 -2540 219 -2537
rect 253 -2542 255 -2524
rect 217 -2563 219 -2560
rect 111 -2566 114 -2564
rect 134 -2566 152 -2564
rect 192 -2566 195 -2564
rect 253 -2565 255 -2562
rect 644 -2574 646 -2546
rect 671 -2558 673 -2546
rect 979 -2558 981 -2555
rect 1006 -2558 1008 -2555
rect 671 -2560 681 -2558
rect 644 -2576 665 -2574
rect 663 -2580 665 -2576
rect -137 -2606 -135 -2602
rect -105 -2606 -103 -2602
rect -338 -2614 -336 -2610
rect -286 -2614 -284 -2610
rect -234 -2614 -232 -2610
rect -182 -2614 -180 -2610
rect 663 -2624 665 -2620
rect 170 -2628 172 -2625
rect 197 -2628 199 -2625
rect -338 -2663 -336 -2654
rect -286 -2663 -284 -2654
rect -234 -2663 -232 -2654
rect -182 -2663 -180 -2654
rect -137 -2666 -135 -2646
rect -105 -2666 -103 -2646
rect -338 -2676 -336 -2672
rect -286 -2676 -284 -2672
rect -234 -2690 -232 -2681
rect -182 -2690 -180 -2681
rect 679 -2637 681 -2560
rect 706 -2576 708 -2573
rect 1309 -2585 1311 -2579
rect 1309 -2587 1329 -2585
rect 706 -2634 708 -2616
rect 979 -2626 981 -2598
rect 1006 -2610 1008 -2598
rect 1309 -2599 1311 -2596
rect 1006 -2612 1016 -2610
rect 979 -2628 1000 -2626
rect 998 -2632 1000 -2628
rect 663 -2639 681 -2637
rect 663 -2645 665 -2639
rect -137 -2690 -135 -2686
rect -105 -2690 -103 -2686
rect 170 -2696 172 -2668
rect 197 -2680 199 -2668
rect 197 -2682 207 -2680
rect 170 -2698 191 -2696
rect 189 -2702 191 -2698
rect -234 -2713 -232 -2710
rect -182 -2713 -180 -2710
rect -338 -2725 -336 -2716
rect -286 -2725 -284 -2716
rect -338 -2737 -336 -2729
rect -286 -2737 -284 -2729
rect -234 -2737 -232 -2729
rect -182 -2737 -180 -2729
rect 189 -2746 191 -2742
rect -338 -2761 -336 -2757
rect -286 -2761 -284 -2757
rect -234 -2761 -232 -2757
rect -182 -2761 -180 -2757
rect 205 -2759 207 -2682
rect 706 -2657 708 -2654
rect 998 -2676 1000 -2672
rect 663 -2688 665 -2685
rect 1014 -2689 1016 -2612
rect 1041 -2628 1043 -2625
rect 1041 -2686 1043 -2668
rect 1309 -2685 1311 -2679
rect 232 -2698 234 -2695
rect 998 -2691 1016 -2689
rect 998 -2697 1000 -2691
rect 1294 -2687 1311 -2685
rect 1294 -2704 1296 -2687
rect 1327 -2704 1329 -2587
rect 1358 -2636 1360 -2633
rect 1358 -2694 1360 -2676
rect 1041 -2709 1043 -2706
rect 1358 -2717 1360 -2714
rect 1294 -2727 1296 -2724
rect 1327 -2727 1329 -2724
rect 232 -2756 234 -2738
rect 998 -2740 1000 -2737
rect 189 -2761 207 -2759
rect 189 -2767 191 -2761
rect 232 -2779 234 -2776
rect 645 -2789 647 -2786
rect 672 -2789 674 -2786
rect 189 -2810 191 -2807
rect 1813 -2813 1815 -2810
rect 645 -2857 647 -2829
rect 672 -2841 674 -2829
rect 980 -2841 982 -2838
rect 1007 -2841 1009 -2838
rect 672 -2843 682 -2841
rect 645 -2859 666 -2857
rect 664 -2863 666 -2859
rect 664 -2907 666 -2903
rect 680 -2920 682 -2843
rect 707 -2859 709 -2856
rect 707 -2917 709 -2899
rect 980 -2909 982 -2881
rect 1007 -2893 1009 -2881
rect 1316 -2888 1318 -2885
rect 1007 -2895 1017 -2893
rect 980 -2911 1001 -2909
rect 999 -2915 1001 -2911
rect 664 -2922 682 -2920
rect 664 -2928 666 -2922
rect 707 -2940 709 -2937
rect 999 -2959 1001 -2955
rect 664 -2971 666 -2968
rect 1015 -2972 1017 -2895
rect 1042 -2911 1044 -2908
rect 1042 -2969 1044 -2951
rect 2287 -2840 2289 -2836
rect 2319 -2840 2321 -2836
rect 2086 -2848 2088 -2844
rect 2138 -2848 2140 -2844
rect 2190 -2848 2192 -2844
rect 2242 -2848 2244 -2844
rect 1813 -2899 1815 -2893
rect 2086 -2897 2088 -2888
rect 2138 -2897 2140 -2888
rect 2190 -2897 2192 -2888
rect 2242 -2897 2244 -2888
rect 1813 -2901 1833 -2899
rect 2287 -2900 2289 -2880
rect 2319 -2900 2321 -2880
rect 1813 -2913 1815 -2910
rect 999 -2974 1017 -2972
rect 999 -2980 1001 -2974
rect 1316 -2974 1318 -2968
rect 1316 -2976 1336 -2974
rect 1316 -2988 1318 -2985
rect 1042 -2992 1044 -2989
rect 999 -3023 1001 -3020
rect 641 -3060 643 -3057
rect 668 -3060 670 -3057
rect 1316 -3074 1318 -3068
rect 1301 -3076 1318 -3074
rect 1301 -3093 1303 -3076
rect 1334 -3093 1336 -2976
rect 1813 -2999 1815 -2993
rect 1798 -3001 1815 -2999
rect 1798 -3018 1800 -3001
rect 1831 -3018 1833 -2901
rect 2086 -2910 2088 -2906
rect 2138 -2910 2140 -2906
rect 1862 -2950 1864 -2947
rect 2190 -2924 2192 -2915
rect 2242 -2924 2244 -2915
rect 2287 -2924 2289 -2920
rect 2319 -2924 2321 -2920
rect 2190 -2947 2192 -2944
rect 2242 -2947 2244 -2944
rect 2086 -2959 2088 -2950
rect 2138 -2959 2140 -2950
rect 2086 -2971 2088 -2963
rect 2138 -2971 2140 -2963
rect 2190 -2971 2192 -2963
rect 2242 -2971 2244 -2963
rect 1862 -3008 1864 -2990
rect 2086 -2995 2088 -2991
rect 2138 -2995 2140 -2991
rect 2190 -2995 2192 -2991
rect 2242 -2995 2244 -2991
rect 1365 -3025 1367 -3022
rect 1862 -3031 1864 -3028
rect 1798 -3041 1800 -3038
rect 1831 -3041 1833 -3038
rect 1608 -3044 1610 -3041
rect 1365 -3083 1367 -3065
rect 641 -3128 643 -3100
rect 668 -3112 670 -3100
rect 668 -3114 678 -3112
rect 1365 -3106 1367 -3103
rect 641 -3130 662 -3128
rect 660 -3134 662 -3130
rect 660 -3178 662 -3174
rect 676 -3191 678 -3114
rect 1301 -3116 1303 -3113
rect 1334 -3116 1336 -3113
rect 703 -3130 705 -3127
rect 1608 -3130 1610 -3124
rect 1608 -3132 1628 -3130
rect 1608 -3144 1610 -3141
rect 703 -3188 705 -3170
rect 660 -3193 678 -3191
rect 660 -3199 662 -3193
rect 703 -3211 705 -3208
rect 1608 -3230 1610 -3224
rect 1593 -3232 1610 -3230
rect 660 -3242 662 -3239
rect 1310 -3243 1312 -3240
rect 1337 -3243 1339 -3240
rect 1593 -3249 1595 -3232
rect 1626 -3249 1628 -3132
rect 1657 -3181 1659 -3178
rect 1657 -3239 1659 -3221
rect 1657 -3262 1659 -3259
rect 1593 -3272 1595 -3269
rect 1626 -3272 1628 -3269
rect 629 -3309 631 -3306
rect 656 -3309 658 -3306
rect 1310 -3311 1312 -3283
rect 1337 -3295 1339 -3283
rect 1337 -3297 1347 -3295
rect 1310 -3313 1331 -3311
rect 1329 -3317 1331 -3313
rect 629 -3377 631 -3349
rect 656 -3361 658 -3349
rect 1329 -3361 1331 -3357
rect 656 -3363 666 -3361
rect 629 -3379 650 -3377
rect 648 -3383 650 -3379
rect 648 -3427 650 -3423
rect 664 -3440 666 -3363
rect 970 -3375 972 -3372
rect 997 -3375 999 -3372
rect 1345 -3374 1347 -3297
rect 1372 -3313 1374 -3310
rect 1372 -3371 1374 -3353
rect 691 -3379 693 -3376
rect 1329 -3376 1347 -3374
rect 1329 -3382 1331 -3376
rect 691 -3437 693 -3419
rect 648 -3442 666 -3440
rect 648 -3448 650 -3442
rect 970 -3443 972 -3415
rect 997 -3427 999 -3415
rect 1372 -3394 1374 -3391
rect 1329 -3425 1331 -3422
rect 997 -3429 1007 -3427
rect 970 -3445 991 -3443
rect 989 -3449 991 -3445
rect 691 -3460 693 -3457
rect 648 -3491 650 -3488
rect 989 -3493 991 -3489
rect 1005 -3506 1007 -3429
rect 1032 -3445 1034 -3442
rect 1032 -3503 1034 -3485
rect 989 -3508 1007 -3506
rect 989 -3514 991 -3508
rect 1032 -3526 1034 -3523
rect 989 -3557 991 -3554
rect 646 -3576 648 -3573
rect 673 -3576 675 -3573
rect 646 -3644 648 -3616
rect 673 -3628 675 -3616
rect 673 -3630 683 -3628
rect 646 -3646 667 -3644
rect 665 -3650 667 -3646
rect 665 -3694 667 -3690
rect 681 -3707 683 -3630
rect 708 -3646 710 -3643
rect 708 -3704 710 -3686
rect 665 -3709 683 -3707
rect 665 -3715 667 -3709
rect 708 -3727 710 -3724
rect 665 -3758 667 -3755
rect 634 -3825 636 -3822
rect 661 -3825 663 -3822
rect 634 -3893 636 -3865
rect 661 -3877 663 -3865
rect 661 -3879 671 -3877
rect 634 -3895 655 -3893
rect 653 -3899 655 -3895
rect 653 -3943 655 -3939
rect 669 -3956 671 -3879
rect 696 -3895 698 -3892
rect 696 -3953 698 -3935
rect 653 -3958 671 -3956
rect 653 -3964 655 -3958
rect 696 -3976 698 -3973
rect 653 -4007 655 -4004
<< polycontact >>
rect 797 1668 802 1673
rect 797 1645 802 1650
rect 797 1623 802 1628
rect 908 1619 913 1624
rect 797 1594 802 1599
rect 999 1603 1004 1608
rect 1064 1613 1069 1618
rect 1173 1619 1178 1624
rect 2845 1641 2850 1646
rect 1049 1510 1054 1515
rect 2845 1618 2850 1623
rect 2845 1596 2850 1601
rect 2956 1592 2961 1597
rect 1235 1564 1240 1569
rect 2845 1567 2850 1572
rect 3047 1576 3052 1581
rect 3112 1586 3117 1591
rect 3221 1592 3226 1597
rect 1192 1553 1197 1558
rect 1113 1509 1118 1514
rect 3097 1483 3102 1488
rect 3283 1537 3288 1542
rect 3240 1526 3245 1531
rect 3161 1482 3166 1487
rect -1528 350 -1523 355
rect -1476 350 -1471 355
rect -1424 350 -1419 355
rect -1372 350 -1367 355
rect -1327 350 -1322 355
rect -1295 350 -1290 355
rect 3767 347 3772 352
rect 3819 347 3824 352
rect 3871 347 3876 352
rect 3923 347 3928 352
rect 3968 347 3973 352
rect -1424 327 -1419 332
rect -1372 327 -1367 332
rect 4000 347 4005 352
rect -1528 288 -1523 293
rect -1476 288 -1471 293
rect 3871 324 3876 329
rect 3923 324 3928 329
rect 3767 285 3772 290
rect 3819 285 3824 290
rect -1528 279 -1523 284
rect -1476 279 -1471 284
rect -1424 279 -1419 284
rect -1372 279 -1367 284
rect 3767 276 3772 281
rect 3819 276 3824 281
rect 3871 276 3876 281
rect 3923 276 3928 281
rect 1419 44 1424 49
rect 1471 44 1476 49
rect 1523 44 1528 49
rect 1575 44 1580 49
rect 1620 44 1625 49
rect 1652 44 1657 49
rect 1056 30 1061 35
rect 1056 7 1061 12
rect 1056 -15 1061 -10
rect 1167 -19 1172 -14
rect -402 -51 -397 -46
rect -350 -51 -345 -46
rect -298 -51 -293 -46
rect -246 -51 -241 -46
rect -201 -51 -196 -46
rect -169 -51 -164 -46
rect 1056 -44 1061 -39
rect 1523 21 1528 26
rect 1575 21 1580 26
rect 1419 -18 1424 -13
rect 1471 -18 1476 -13
rect 1419 -27 1424 -22
rect 1471 -27 1476 -22
rect 1523 -27 1528 -22
rect 1575 -27 1580 -22
rect -298 -74 -293 -69
rect -246 -74 -241 -69
rect -402 -113 -397 -108
rect -350 -113 -345 -108
rect -402 -122 -397 -117
rect -350 -122 -345 -117
rect -298 -122 -293 -117
rect -246 -122 -241 -117
rect 143 -169 148 -164
rect 143 -192 148 -187
rect 816 -148 821 -143
rect 143 -214 148 -209
rect 254 -218 259 -213
rect 143 -243 148 -238
rect 446 -215 451 -210
rect 801 -251 806 -246
rect 508 -270 513 -265
rect 1051 -190 1056 -185
rect 1051 -213 1056 -208
rect 1051 -235 1056 -230
rect 865 -252 870 -247
rect 1162 -239 1167 -234
rect 465 -281 470 -276
rect -406 -306 -401 -301
rect -354 -306 -349 -301
rect -302 -306 -297 -301
rect -250 -306 -245 -301
rect -205 -306 -200 -301
rect -173 -306 -168 -301
rect -302 -329 -297 -324
rect -250 -329 -245 -324
rect 1051 -264 1056 -259
rect 1434 -232 1439 -227
rect 1486 -232 1491 -227
rect 1538 -232 1543 -227
rect 1590 -232 1595 -227
rect 1635 -232 1640 -227
rect 1667 -232 1672 -227
rect 1538 -255 1543 -250
rect 1590 -255 1595 -250
rect 1434 -294 1439 -289
rect 1486 -294 1491 -289
rect 1434 -303 1439 -298
rect 1486 -303 1491 -298
rect 1538 -303 1543 -298
rect 1590 -303 1595 -298
rect -406 -368 -401 -363
rect -354 -368 -349 -363
rect -406 -377 -401 -372
rect -354 -377 -349 -372
rect -302 -377 -297 -372
rect -250 -377 -245 -372
rect 171 -377 176 -372
rect 233 -432 238 -427
rect 190 -443 195 -438
rect 960 -795 965 -790
rect 626 -866 631 -861
rect -309 -888 -304 -883
rect -257 -888 -252 -883
rect -205 -888 -200 -883
rect -153 -888 -148 -883
rect -108 -888 -103 -883
rect -76 -888 -71 -883
rect -205 -911 -200 -906
rect -153 -911 -148 -906
rect 945 -898 950 -893
rect 688 -921 693 -916
rect 1211 -797 1216 -792
rect 1009 -899 1014 -894
rect 1196 -900 1201 -895
rect 645 -932 650 -927
rect -309 -950 -304 -945
rect -257 -950 -252 -945
rect -309 -959 -304 -954
rect -257 -959 -252 -954
rect -205 -959 -200 -954
rect -153 -959 -148 -954
rect 131 -955 136 -950
rect 131 -978 136 -973
rect 1260 -901 1265 -896
rect 1818 -905 1823 -900
rect 1870 -905 1875 -900
rect 1922 -905 1927 -900
rect 1974 -905 1979 -900
rect 2019 -905 2024 -900
rect 2051 -905 2056 -900
rect 1503 -920 1508 -915
rect 1503 -943 1508 -938
rect 1503 -965 1508 -960
rect 1614 -969 1619 -964
rect 131 -1000 136 -995
rect 242 -1004 247 -999
rect 131 -1029 136 -1024
rect 1503 -994 1508 -989
rect 1922 -928 1927 -923
rect 1974 -928 1979 -923
rect 1818 -967 1823 -962
rect 1870 -967 1875 -962
rect 1818 -976 1823 -971
rect 1870 -976 1875 -971
rect 1922 -976 1927 -971
rect 1974 -976 1979 -971
rect -328 -1111 -323 -1106
rect -276 -1111 -271 -1106
rect -224 -1111 -219 -1106
rect -172 -1111 -167 -1106
rect -127 -1111 -122 -1106
rect -95 -1111 -90 -1106
rect -3556 -1189 -3551 -1184
rect -3556 -1212 -3551 -1207
rect -3556 -1234 -3551 -1229
rect -3445 -1238 -3440 -1233
rect -3556 -1263 -3551 -1258
rect -224 -1134 -219 -1129
rect -172 -1134 -167 -1129
rect 549 -1111 554 -1106
rect 159 -1163 164 -1158
rect -328 -1173 -323 -1168
rect -276 -1173 -271 -1168
rect -328 -1182 -323 -1177
rect -276 -1182 -271 -1177
rect -224 -1182 -219 -1177
rect -172 -1182 -167 -1177
rect -3354 -1254 -3349 -1249
rect -3289 -1244 -3284 -1239
rect -3180 -1238 -3175 -1233
rect -3304 -1347 -3299 -1342
rect 767 -1111 772 -1106
rect 611 -1166 616 -1161
rect 568 -1177 573 -1172
rect 221 -1218 226 -1213
rect 829 -1166 834 -1161
rect 786 -1177 791 -1172
rect 178 -1229 183 -1224
rect -3118 -1293 -3113 -1288
rect -3161 -1304 -3156 -1299
rect -3240 -1348 -3235 -1343
rect 561 -1426 566 -1421
rect -328 -1449 -323 -1444
rect -276 -1449 -271 -1444
rect -224 -1449 -219 -1444
rect -172 -1449 -167 -1444
rect -127 -1449 -122 -1444
rect -95 -1449 -90 -1444
rect -224 -1472 -219 -1467
rect -172 -1472 -167 -1467
rect 623 -1481 628 -1476
rect 580 -1492 585 -1487
rect -328 -1511 -323 -1506
rect -276 -1511 -271 -1506
rect -328 -1520 -323 -1515
rect -276 -1520 -271 -1515
rect -224 -1520 -219 -1515
rect -172 -1520 -167 -1515
rect 1080 -1520 1085 -1515
rect 140 -1615 145 -1610
rect 140 -1638 145 -1633
rect 1065 -1623 1070 -1618
rect 140 -1660 145 -1655
rect 251 -1664 256 -1659
rect 140 -1689 145 -1684
rect 798 -1656 803 -1651
rect 1129 -1624 1134 -1619
rect 562 -1709 567 -1704
rect -343 -1786 -338 -1781
rect -291 -1786 -286 -1781
rect -239 -1786 -234 -1781
rect -187 -1786 -182 -1781
rect -142 -1786 -137 -1781
rect -110 -1786 -105 -1781
rect -239 -1809 -234 -1804
rect -187 -1809 -182 -1804
rect 1684 -1656 1689 -1651
rect 1377 -1673 1382 -1668
rect 860 -1711 865 -1706
rect 817 -1722 822 -1717
rect 624 -1764 629 -1759
rect 581 -1775 586 -1770
rect 168 -1823 173 -1818
rect -343 -1848 -338 -1843
rect -291 -1848 -286 -1843
rect -343 -1857 -338 -1852
rect -291 -1857 -286 -1852
rect -239 -1857 -234 -1852
rect -187 -1857 -182 -1852
rect 1362 -1776 1367 -1771
rect 1684 -1679 1689 -1674
rect 2007 -1655 2012 -1650
rect 2059 -1655 2064 -1650
rect 2111 -1655 2116 -1650
rect 2163 -1655 2168 -1650
rect 2208 -1655 2213 -1650
rect 2240 -1655 2245 -1650
rect 1684 -1701 1689 -1696
rect 1795 -1705 1800 -1700
rect 1684 -1730 1689 -1725
rect 2111 -1678 2116 -1673
rect 2163 -1678 2168 -1673
rect 2007 -1717 2012 -1712
rect 2059 -1717 2064 -1712
rect 2007 -1726 2012 -1721
rect 2059 -1726 2064 -1721
rect 2111 -1726 2116 -1721
rect 2163 -1726 2168 -1721
rect 1426 -1777 1431 -1772
rect 1091 -1820 1096 -1815
rect 230 -1878 235 -1873
rect 807 -1867 812 -1862
rect 187 -1889 192 -1884
rect 869 -1922 874 -1917
rect 1076 -1923 1081 -1918
rect 826 -1933 831 -1928
rect 558 -1980 563 -1975
rect 1140 -1924 1145 -1919
rect 620 -2035 625 -2030
rect 577 -2046 582 -2041
rect 546 -2229 551 -2224
rect 608 -2284 613 -2279
rect 565 -2295 570 -2290
rect -343 -2393 -338 -2388
rect -291 -2393 -286 -2388
rect -239 -2393 -234 -2388
rect -187 -2393 -182 -2388
rect -142 -2393 -137 -2388
rect -110 -2393 -105 -2388
rect -239 -2416 -234 -2411
rect -187 -2416 -182 -2411
rect -343 -2455 -338 -2450
rect -291 -2455 -286 -2450
rect -343 -2464 -338 -2459
rect -291 -2464 -286 -2459
rect -239 -2464 -234 -2459
rect -187 -2464 -182 -2459
rect 137 -2490 142 -2485
rect 137 -2513 142 -2508
rect 137 -2535 142 -2530
rect 248 -2539 253 -2534
rect 137 -2564 142 -2559
rect 639 -2576 644 -2571
rect -343 -2663 -338 -2658
rect -291 -2663 -286 -2658
rect -239 -2663 -234 -2658
rect -187 -2663 -182 -2658
rect -142 -2663 -137 -2658
rect -110 -2663 -105 -2658
rect -239 -2686 -234 -2681
rect -187 -2686 -182 -2681
rect 1304 -2587 1309 -2582
rect 701 -2631 706 -2626
rect 974 -2628 979 -2623
rect 658 -2642 663 -2637
rect 165 -2698 170 -2693
rect -343 -2725 -338 -2720
rect -291 -2725 -286 -2720
rect -343 -2734 -338 -2729
rect -291 -2734 -286 -2729
rect -239 -2734 -234 -2729
rect -187 -2734 -182 -2729
rect 1036 -2683 1041 -2678
rect 993 -2694 998 -2689
rect 1289 -2690 1294 -2685
rect 1353 -2691 1358 -2686
rect 227 -2753 232 -2748
rect 184 -2764 189 -2759
rect 640 -2859 645 -2854
rect 702 -2914 707 -2909
rect 975 -2911 980 -2906
rect 659 -2925 664 -2920
rect 1037 -2966 1042 -2961
rect 1808 -2901 1813 -2896
rect 2081 -2897 2086 -2892
rect 2133 -2897 2138 -2892
rect 2185 -2897 2190 -2892
rect 2237 -2897 2242 -2892
rect 2282 -2897 2287 -2892
rect 2314 -2897 2319 -2892
rect 994 -2977 999 -2972
rect 1311 -2976 1316 -2971
rect 1296 -3079 1301 -3074
rect 1793 -3004 1798 -2999
rect 2185 -2920 2190 -2915
rect 2237 -2920 2242 -2915
rect 2081 -2959 2086 -2954
rect 2133 -2959 2138 -2954
rect 2081 -2968 2086 -2963
rect 2133 -2968 2138 -2963
rect 2185 -2968 2190 -2963
rect 2237 -2968 2242 -2963
rect 1857 -3005 1862 -3000
rect 1360 -3080 1365 -3075
rect 636 -3130 641 -3125
rect 1603 -3132 1608 -3127
rect 698 -3185 703 -3180
rect 655 -3196 660 -3191
rect 1588 -3235 1593 -3230
rect 1652 -3236 1657 -3231
rect 1305 -3313 1310 -3308
rect 624 -3379 629 -3374
rect 1367 -3368 1372 -3363
rect 1324 -3379 1329 -3374
rect 686 -3434 691 -3429
rect 643 -3445 648 -3440
rect 965 -3445 970 -3440
rect 1027 -3500 1032 -3495
rect 984 -3511 989 -3506
rect 641 -3646 646 -3641
rect 703 -3701 708 -3696
rect 660 -3712 665 -3707
rect 629 -3895 634 -3890
rect 691 -3950 696 -3945
rect 648 -3961 653 -3956
<< metal1 >>
rect 1056 1712 1083 1715
rect 1056 1708 1059 1712
rect 1063 1708 1076 1712
rect 1080 1708 1083 1712
rect 1056 1706 1083 1708
rect 1064 1701 1068 1706
rect 900 1685 927 1688
rect 900 1681 903 1685
rect 907 1681 920 1685
rect 924 1681 927 1685
rect 900 1679 927 1681
rect 908 1674 912 1679
rect 797 1666 802 1668
rect 762 1661 802 1666
rect 762 1657 768 1658
rect 762 1653 763 1657
rect 767 1653 768 1657
rect 762 1650 768 1653
rect 797 1650 802 1661
rect 857 1655 866 1658
rect 857 1651 859 1655
rect 863 1651 866 1655
rect 880 1651 893 1654
rect 857 1650 866 1651
rect 762 1646 774 1650
rect 762 1636 768 1646
rect 852 1646 866 1650
rect 794 1638 812 1642
rect 857 1638 866 1646
rect 762 1632 763 1636
rect 767 1632 768 1636
rect 762 1631 768 1632
rect 797 1628 802 1638
rect 857 1634 859 1638
rect 863 1634 866 1638
rect 857 1631 866 1634
rect 872 1628 876 1631
rect 826 1624 876 1628
rect 826 1619 830 1624
rect 762 1614 830 1619
rect 880 1618 884 1631
rect 887 1624 893 1651
rect 991 1669 1018 1672
rect 991 1665 994 1669
rect 998 1665 1011 1669
rect 1015 1665 1018 1669
rect 991 1663 1018 1665
rect 916 1624 920 1634
rect 999 1658 1003 1663
rect 887 1619 908 1624
rect 916 1619 927 1624
rect 762 1606 768 1607
rect 762 1602 763 1606
rect 767 1602 768 1606
rect 762 1599 768 1602
rect 797 1599 802 1614
rect 857 1604 866 1607
rect 857 1600 859 1604
rect 863 1600 866 1604
rect 857 1599 866 1600
rect 762 1595 774 1599
rect 762 1585 768 1595
rect 852 1595 866 1599
rect 794 1587 812 1591
rect 857 1587 866 1595
rect 762 1581 763 1585
rect 767 1581 768 1585
rect 762 1580 768 1581
rect 797 1567 802 1587
rect 857 1583 859 1587
rect 863 1583 866 1587
rect 857 1580 866 1583
rect 916 1616 920 1619
rect 1165 1700 1219 1703
rect 1165 1696 1168 1700
rect 1172 1696 1185 1700
rect 1189 1696 1195 1700
rect 1199 1696 1212 1700
rect 1216 1696 1219 1700
rect 1165 1694 1219 1696
rect 1173 1689 1177 1694
rect 1200 1689 1204 1694
rect 3104 1685 3131 1688
rect 3104 1681 3107 1685
rect 3111 1681 3124 1685
rect 3128 1681 3131 1685
rect 3104 1679 3131 1681
rect 3112 1674 3116 1679
rect 2948 1658 2975 1661
rect 2948 1654 2951 1658
rect 2955 1654 2968 1658
rect 2972 1654 2975 1658
rect 2948 1652 2975 1654
rect 1181 1629 1185 1649
rect 1208 1629 1212 1649
rect 2956 1647 2960 1652
rect 2845 1639 2850 1641
rect 2810 1634 2850 1639
rect 1227 1630 1254 1633
rect 1181 1625 1222 1629
rect 872 1567 876 1598
rect 1007 1608 1011 1618
rect 1047 1613 1064 1618
rect 1072 1609 1076 1621
rect 1166 1619 1173 1624
rect 1200 1615 1204 1625
rect 991 1603 999 1608
rect 1007 1603 1020 1608
rect 1064 1605 1076 1609
rect 1007 1600 1011 1603
rect 908 1590 912 1596
rect 900 1589 927 1590
rect 900 1585 901 1589
rect 905 1585 922 1589
rect 926 1585 927 1589
rect 900 1584 927 1585
rect 1064 1601 1068 1605
rect 999 1574 1003 1580
rect 991 1573 1018 1574
rect 991 1569 992 1573
rect 996 1569 1013 1573
rect 1017 1569 1018 1573
rect 991 1568 1018 1569
rect 797 1564 876 1567
rect 1105 1575 1132 1578
rect 1105 1571 1108 1575
rect 1112 1571 1125 1575
rect 1129 1571 1132 1575
rect 1105 1569 1132 1571
rect 1192 1569 1196 1575
rect 1217 1569 1222 1625
rect 1227 1626 1230 1630
rect 1234 1626 1247 1630
rect 1251 1626 1254 1630
rect 1227 1624 1254 1626
rect 2810 1630 2816 1631
rect 2810 1626 2811 1630
rect 2815 1626 2816 1630
rect 1235 1619 1239 1624
rect 2810 1623 2816 1626
rect 2845 1623 2850 1634
rect 2905 1628 2914 1631
rect 2905 1624 2907 1628
rect 2911 1624 2914 1628
rect 2928 1624 2941 1627
rect 2905 1623 2914 1624
rect 2810 1619 2822 1623
rect 2810 1609 2816 1619
rect 2900 1619 2914 1623
rect 2842 1611 2860 1615
rect 2905 1611 2914 1619
rect 2810 1605 2811 1609
rect 2815 1605 2816 1609
rect 2810 1604 2816 1605
rect 2845 1601 2850 1611
rect 2905 1607 2907 1611
rect 2911 1607 2914 1611
rect 2905 1604 2914 1607
rect 2920 1601 2924 1604
rect 2874 1597 2924 1601
rect 2874 1592 2878 1597
rect 2810 1587 2878 1592
rect 2928 1591 2932 1604
rect 2935 1597 2941 1624
rect 3039 1642 3066 1645
rect 3039 1638 3042 1642
rect 3046 1638 3059 1642
rect 3063 1638 3066 1642
rect 3039 1636 3066 1638
rect 2964 1597 2968 1607
rect 3047 1631 3051 1636
rect 2935 1592 2956 1597
rect 2964 1592 2975 1597
rect 1243 1569 1247 1579
rect 2810 1579 2816 1580
rect 2810 1575 2811 1579
rect 2815 1575 2816 1579
rect 2810 1572 2816 1575
rect 2845 1572 2850 1587
rect 2905 1577 2914 1580
rect 2905 1573 2907 1577
rect 2911 1573 2914 1577
rect 2905 1572 2914 1573
rect 1113 1564 1117 1569
rect 1192 1565 1206 1569
rect 1200 1564 1206 1565
rect 1217 1564 1235 1569
rect 1243 1564 1256 1569
rect 2810 1568 2822 1572
rect 1166 1553 1192 1558
rect 1200 1550 1204 1564
rect 1243 1561 1247 1564
rect 1040 1510 1049 1515
rect 1072 1514 1076 1521
rect 1121 1514 1125 1524
rect 1072 1509 1113 1514
rect 1121 1509 1132 1514
rect 2810 1558 2816 1568
rect 2900 1568 2914 1572
rect 2842 1560 2860 1564
rect 2905 1560 2914 1568
rect 2810 1554 2811 1558
rect 2815 1554 2816 1558
rect 2810 1553 2816 1554
rect 1235 1535 1239 1541
rect 2845 1540 2850 1560
rect 2905 1556 2907 1560
rect 2911 1556 2914 1560
rect 2905 1553 2914 1556
rect 2964 1589 2968 1592
rect 3213 1673 3267 1676
rect 3213 1669 3216 1673
rect 3220 1669 3233 1673
rect 3237 1669 3243 1673
rect 3247 1669 3260 1673
rect 3264 1669 3267 1673
rect 3213 1667 3267 1669
rect 3221 1662 3225 1667
rect 3248 1662 3252 1667
rect 3229 1602 3233 1622
rect 3256 1602 3260 1622
rect 3275 1603 3302 1606
rect 3229 1598 3270 1602
rect 2920 1540 2924 1571
rect 3055 1581 3059 1591
rect 3095 1586 3112 1591
rect 3120 1582 3124 1594
rect 3214 1592 3221 1597
rect 3248 1588 3252 1598
rect 3039 1576 3047 1581
rect 3055 1576 3068 1581
rect 3112 1578 3124 1582
rect 3055 1573 3059 1576
rect 2956 1563 2960 1569
rect 2948 1562 2975 1563
rect 2948 1558 2949 1562
rect 2953 1558 2970 1562
rect 2974 1558 2975 1562
rect 2948 1557 2975 1558
rect 3112 1574 3116 1578
rect 3047 1547 3051 1553
rect 3039 1546 3066 1547
rect 3039 1542 3040 1546
rect 3044 1542 3061 1546
rect 3065 1542 3066 1546
rect 3039 1541 3066 1542
rect 2845 1537 2924 1540
rect 1227 1534 1254 1535
rect 1227 1530 1228 1534
rect 1232 1530 1249 1534
rect 1253 1530 1254 1534
rect 1227 1529 1254 1530
rect 1072 1506 1076 1509
rect 1121 1506 1125 1509
rect 1057 1502 1094 1506
rect 1057 1496 1061 1502
rect 1090 1496 1094 1502
rect 1192 1504 1196 1510
rect 1184 1503 1211 1504
rect 1184 1499 1185 1503
rect 1189 1499 1206 1503
rect 1210 1499 1211 1503
rect 1184 1498 1211 1499
rect 3153 1548 3180 1551
rect 3153 1544 3156 1548
rect 3160 1544 3173 1548
rect 3177 1544 3180 1548
rect 3153 1542 3180 1544
rect 3240 1542 3244 1548
rect 3265 1542 3270 1598
rect 3275 1599 3278 1603
rect 3282 1599 3295 1603
rect 3299 1599 3302 1603
rect 3275 1597 3302 1599
rect 3283 1592 3287 1597
rect 3291 1542 3295 1552
rect 3161 1537 3165 1542
rect 3240 1538 3254 1542
rect 3248 1537 3254 1538
rect 3265 1537 3283 1542
rect 3291 1537 3304 1542
rect 3214 1526 3240 1531
rect 3248 1523 3252 1537
rect 3291 1534 3295 1537
rect 1113 1480 1117 1486
rect 3088 1483 3097 1488
rect 3120 1487 3124 1494
rect 3169 1487 3173 1497
rect 3120 1482 3161 1487
rect 3169 1482 3180 1487
rect 3283 1508 3287 1514
rect 3275 1507 3302 1508
rect 3275 1503 3276 1507
rect 3280 1503 3297 1507
rect 3301 1503 3302 1507
rect 3275 1502 3302 1503
rect 1105 1479 1132 1480
rect 3120 1479 3124 1482
rect 3169 1479 3173 1482
rect 1049 1470 1053 1476
rect 1082 1470 1086 1476
rect 1105 1475 1106 1479
rect 1110 1475 1127 1479
rect 1131 1475 1132 1479
rect 1105 1474 1132 1475
rect 3105 1475 3142 1479
rect 1041 1469 1068 1470
rect 1041 1465 1042 1469
rect 1046 1465 1063 1469
rect 1067 1465 1068 1469
rect 1041 1464 1068 1465
rect 1074 1469 1101 1470
rect 3105 1469 3109 1475
rect 3138 1469 3142 1475
rect 1074 1465 1075 1469
rect 1079 1465 1096 1469
rect 1100 1465 1101 1469
rect 1074 1464 1101 1465
rect 3240 1477 3244 1483
rect 3232 1476 3259 1477
rect 3232 1472 3233 1476
rect 3237 1472 3254 1476
rect 3258 1472 3259 1476
rect 3232 1471 3259 1472
rect 3161 1453 3165 1459
rect 3153 1452 3180 1453
rect 3097 1443 3101 1449
rect 3130 1443 3134 1449
rect 3153 1448 3154 1452
rect 3158 1448 3175 1452
rect 3179 1448 3180 1452
rect 3153 1447 3180 1448
rect 3089 1442 3116 1443
rect 3089 1438 3090 1442
rect 3094 1438 3111 1442
rect 3115 1438 3116 1442
rect 3089 1437 3116 1438
rect 3122 1442 3149 1443
rect 3122 1438 3123 1442
rect 3127 1438 3144 1442
rect 3148 1438 3149 1442
rect 3122 1437 3149 1438
rect -1337 419 -1273 422
rect -1337 415 -1334 419
rect -1330 415 -1312 419
rect -1308 415 -1302 419
rect -1298 415 -1280 419
rect -1276 415 -1273 419
rect -1538 411 -1350 414
rect -1337 413 -1273 415
rect 3958 416 4022 419
rect -1538 407 -1535 411
rect -1531 407 -1513 411
rect -1509 407 -1483 411
rect -1479 407 -1461 411
rect -1457 407 -1431 411
rect -1427 407 -1409 411
rect -1405 407 -1379 411
rect -1375 407 -1357 411
rect -1353 407 -1350 411
rect -1538 405 -1350 407
rect -1327 407 -1323 413
rect -1295 407 -1291 413
rect 3958 412 3961 416
rect 3965 412 3983 416
rect 3987 412 3993 416
rect 3997 412 4015 416
rect 4019 412 4022 416
rect 3757 408 3945 411
rect 3958 410 4022 412
rect -1528 399 -1524 405
rect -1476 399 -1472 405
rect -1424 399 -1420 405
rect -1372 399 -1368 405
rect 3757 404 3760 408
rect 3764 404 3782 408
rect 3786 404 3812 408
rect 3816 404 3834 408
rect 3838 404 3864 408
rect 3868 404 3886 408
rect 3890 404 3916 408
rect 3920 404 3938 408
rect 3942 404 3945 408
rect 3757 402 3945 404
rect 3968 404 3972 410
rect 4000 404 4004 410
rect -1551 350 -1528 355
rect -1551 284 -1546 350
rect -1520 346 -1516 359
rect -1528 342 -1516 346
rect -1498 350 -1476 355
rect -1528 337 -1524 342
rect -1533 288 -1528 293
rect -1520 284 -1516 297
rect -1498 284 -1493 350
rect -1468 346 -1464 359
rect -1416 355 -1412 359
rect -1364 355 -1360 359
rect -1319 355 -1315 367
rect -1287 355 -1283 367
rect 3767 396 3771 402
rect 3819 396 3823 402
rect 3871 396 3875 402
rect 3923 396 3927 402
rect -1476 342 -1464 346
rect -1446 350 -1424 355
rect -1416 350 -1372 355
rect -1364 350 -1327 355
rect -1319 350 -1295 355
rect -1287 350 -1273 355
rect -1476 337 -1472 342
rect -1481 288 -1476 293
rect -1468 284 -1464 297
rect -1446 284 -1441 350
rect -1427 327 -1424 332
rect -1416 323 -1412 350
rect -1424 292 -1420 303
rect -1424 288 -1412 292
rect -1551 279 -1528 284
rect -1520 279 -1476 284
rect -1468 279 -1424 284
rect -1520 276 -1516 279
rect -1468 276 -1464 279
rect -1416 276 -1412 288
rect -1394 284 -1389 350
rect -1375 327 -1372 332
rect -1364 323 -1360 350
rect -1319 347 -1315 350
rect -1287 347 -1283 350
rect 3744 347 3767 352
rect -1327 320 -1323 327
rect -1295 320 -1291 327
rect -1337 318 -1273 320
rect -1337 314 -1335 318
rect -1331 314 -1311 318
rect -1307 314 -1303 318
rect -1299 314 -1279 318
rect -1275 314 -1273 318
rect -1337 312 -1273 314
rect -1372 292 -1368 303
rect -1372 288 -1360 292
rect -1394 279 -1372 284
rect -1364 276 -1360 288
rect 3744 281 3749 347
rect 3775 343 3779 356
rect 3767 339 3779 343
rect 3797 347 3819 352
rect 3767 334 3771 339
rect 3762 285 3767 290
rect 3775 281 3779 294
rect 3797 281 3802 347
rect 3827 343 3831 356
rect 3879 352 3883 356
rect 3931 352 3935 356
rect 3976 352 3980 364
rect 4008 352 4012 364
rect 3819 339 3831 343
rect 3849 347 3871 352
rect 3879 347 3923 352
rect 3931 347 3968 352
rect 3976 347 4000 352
rect 4008 347 4022 352
rect 3819 334 3823 339
rect 3814 285 3819 290
rect 3827 281 3831 294
rect 3849 281 3854 347
rect 3868 324 3871 329
rect 3879 320 3883 347
rect 3871 289 3875 300
rect 3871 285 3883 289
rect 3744 276 3767 281
rect 3775 276 3819 281
rect 3827 276 3871 281
rect 3775 273 3779 276
rect 3827 273 3831 276
rect 3879 273 3883 285
rect 3901 281 3906 347
rect 3920 324 3923 329
rect 3931 320 3935 347
rect 3976 344 3980 347
rect 4008 344 4012 347
rect 3968 317 3972 324
rect 4000 317 4004 324
rect 3958 315 4022 317
rect 3958 311 3960 315
rect 3964 311 3984 315
rect 3988 311 3992 315
rect 3996 311 4016 315
rect 4020 311 4022 315
rect 3958 309 4022 311
rect 3923 289 3927 300
rect 3923 285 3935 289
rect 3901 276 3923 281
rect 3931 273 3935 285
rect -1528 248 -1524 256
rect -1476 248 -1472 256
rect -1424 248 -1420 256
rect -1372 248 -1368 256
rect -1538 247 -1350 248
rect -1538 243 -1511 247
rect -1507 243 -1459 247
rect -1455 243 -1407 247
rect -1403 243 -1355 247
rect -1351 243 -1350 247
rect 3767 245 3771 253
rect 3819 245 3823 253
rect 3871 245 3875 253
rect 3923 245 3927 253
rect -1538 242 -1350 243
rect 3757 244 3945 245
rect 3757 240 3784 244
rect 3788 240 3836 244
rect 3840 240 3888 244
rect 3892 240 3940 244
rect 3944 240 3945 244
rect 3757 239 3945 240
rect -1545 229 -1538 234
rect -1533 229 -1486 234
rect -1481 229 -1432 234
rect -1427 229 -1380 234
rect 3750 226 3757 231
rect 3762 226 3809 231
rect 3814 226 3863 231
rect 3868 226 3915 231
rect 1610 113 1674 116
rect 1610 109 1613 113
rect 1617 109 1635 113
rect 1639 109 1645 113
rect 1649 109 1667 113
rect 1671 109 1674 113
rect 1409 105 1597 108
rect 1610 107 1674 109
rect 1409 101 1412 105
rect 1416 101 1434 105
rect 1438 101 1464 105
rect 1468 101 1486 105
rect 1490 101 1516 105
rect 1520 101 1538 105
rect 1542 101 1568 105
rect 1572 101 1590 105
rect 1594 101 1597 105
rect 1409 99 1597 101
rect 1620 101 1624 107
rect 1652 101 1656 107
rect 1419 93 1423 99
rect 1471 93 1475 99
rect 1523 93 1527 99
rect 1575 93 1579 99
rect 1159 47 1186 50
rect 1159 43 1162 47
rect 1166 43 1179 47
rect 1183 43 1186 47
rect 1159 41 1186 43
rect 1396 44 1419 49
rect 1167 36 1171 41
rect 429 31 936 33
rect -31 26 299 30
rect 413 30 936 31
rect 304 29 936 30
rect 304 26 440 29
rect 458 28 936 29
rect 1056 28 1061 30
rect 413 25 440 26
rect 926 23 1061 28
rect -211 18 -147 21
rect -211 14 -208 18
rect -204 14 -186 18
rect -182 14 -176 18
rect -172 14 -154 18
rect -150 14 -147 18
rect -412 10 -224 13
rect -211 12 -147 14
rect 1021 19 1027 20
rect 1021 15 1022 19
rect 1026 15 1027 19
rect 1021 12 1027 15
rect 1056 12 1061 23
rect 1116 17 1125 20
rect 1116 13 1118 17
rect 1122 13 1125 17
rect 1139 13 1152 16
rect 1116 12 1125 13
rect -412 6 -409 10
rect -405 6 -387 10
rect -383 6 -357 10
rect -353 6 -335 10
rect -331 6 -305 10
rect -301 6 -283 10
rect -279 6 -253 10
rect -249 6 -231 10
rect -227 6 -224 10
rect -412 4 -224 6
rect -201 6 -197 12
rect -169 6 -165 12
rect 1021 8 1033 12
rect -402 -2 -398 4
rect -350 -2 -346 4
rect -298 -2 -294 4
rect -246 -2 -242 4
rect 1021 -2 1027 8
rect 1111 8 1125 12
rect 1053 0 1071 4
rect 1116 0 1125 8
rect 1021 -6 1022 -2
rect 1026 -6 1027 -2
rect 1021 -7 1027 -6
rect 1056 -10 1061 0
rect 1116 -4 1118 0
rect 1122 -4 1125 0
rect 1116 -7 1125 -4
rect 1131 -10 1135 -7
rect 429 -17 936 -14
rect 1085 -14 1135 -10
rect 313 -19 936 -17
rect 1085 -19 1089 -14
rect 313 -22 438 -19
rect 411 -23 438 -22
rect 926 -24 1089 -19
rect 1139 -20 1143 -7
rect 1146 -14 1152 13
rect 1175 -14 1179 -4
rect 1396 -14 1401 44
rect 1427 40 1431 53
rect 1419 36 1431 40
rect 1449 44 1471 49
rect 1419 31 1423 36
rect 1146 -19 1167 -14
rect 1175 -19 1401 -14
rect 1414 -18 1419 -13
rect -425 -51 -402 -46
rect -425 -117 -420 -51
rect -394 -55 -390 -42
rect -402 -59 -390 -55
rect -372 -51 -350 -46
rect -402 -64 -398 -59
rect -407 -113 -402 -108
rect -394 -117 -390 -104
rect -372 -117 -367 -51
rect -342 -55 -338 -42
rect -290 -46 -286 -42
rect -238 -46 -234 -42
rect -193 -46 -189 -34
rect -161 -46 -157 -34
rect 1021 -32 1027 -31
rect 1021 -36 1022 -32
rect 1026 -36 1027 -32
rect 1021 -39 1027 -36
rect 1056 -39 1061 -24
rect 1116 -34 1125 -31
rect 1116 -38 1118 -34
rect 1122 -38 1125 -34
rect 1116 -39 1125 -38
rect 1021 -43 1033 -39
rect -350 -59 -338 -55
rect -320 -51 -298 -46
rect -290 -51 -246 -46
rect -238 -51 -201 -46
rect -193 -51 -169 -46
rect -161 -51 -9 -46
rect -350 -64 -346 -59
rect -355 -113 -350 -108
rect -342 -117 -338 -104
rect -320 -117 -315 -51
rect -301 -74 -298 -69
rect -290 -78 -286 -51
rect -298 -109 -294 -98
rect -298 -113 -286 -109
rect -425 -122 -402 -117
rect -394 -122 -350 -117
rect -342 -122 -298 -117
rect -394 -125 -390 -122
rect -342 -125 -338 -122
rect -290 -125 -286 -113
rect -268 -117 -263 -51
rect -249 -74 -246 -69
rect -238 -78 -234 -51
rect -193 -54 -189 -51
rect -161 -54 -157 -51
rect -147 -52 -9 -51
rect -201 -81 -197 -74
rect -169 -81 -165 -74
rect -211 -83 -147 -81
rect -211 -87 -209 -83
rect -205 -87 -185 -83
rect -181 -87 -177 -83
rect -173 -87 -153 -83
rect -149 -87 -147 -83
rect -211 -89 -147 -87
rect -246 -109 -242 -98
rect -246 -113 -234 -109
rect -268 -122 -246 -117
rect -238 -125 -234 -113
rect -402 -153 -398 -145
rect -350 -153 -346 -145
rect -298 -153 -294 -145
rect -246 -153 -242 -145
rect -412 -154 -224 -153
rect -412 -158 -385 -154
rect -381 -158 -333 -154
rect -329 -158 -281 -154
rect -277 -158 -229 -154
rect -225 -158 -224 -154
rect -412 -159 -224 -158
rect -419 -172 -412 -167
rect -407 -172 -360 -167
rect -355 -172 -306 -167
rect -301 -172 -254 -167
rect -19 -171 -9 -52
rect 808 -49 835 -46
rect 808 -53 811 -49
rect 815 -53 828 -49
rect 832 -53 835 -49
rect 808 -55 835 -53
rect 1021 -53 1027 -43
rect 1111 -43 1125 -39
rect 1053 -51 1071 -47
rect 1116 -51 1125 -43
rect 816 -60 820 -55
rect 1021 -57 1022 -53
rect 1026 -57 1027 -53
rect 1021 -58 1027 -57
rect 438 -134 492 -131
rect 438 -138 441 -134
rect 445 -138 458 -134
rect 462 -138 468 -134
rect 472 -138 485 -134
rect 489 -138 492 -134
rect 438 -140 492 -138
rect 1056 -71 1061 -51
rect 1116 -55 1118 -51
rect 1122 -55 1125 -51
rect 1116 -58 1125 -55
rect 1175 -22 1179 -19
rect 1221 -21 1401 -19
rect 1131 -71 1135 -40
rect 1396 -22 1401 -21
rect 1427 -22 1431 -9
rect 1449 -22 1454 44
rect 1479 40 1483 53
rect 1531 49 1535 53
rect 1583 49 1587 53
rect 1628 49 1632 61
rect 1660 49 1664 61
rect 1471 36 1483 40
rect 1501 44 1523 49
rect 1531 44 1575 49
rect 1583 44 1620 49
rect 1628 44 1652 49
rect 1660 44 1674 49
rect 1471 31 1475 36
rect 1466 -18 1471 -13
rect 1479 -22 1483 -9
rect 1501 -22 1506 44
rect 1520 21 1523 26
rect 1531 17 1535 44
rect 1523 -14 1527 -3
rect 1523 -18 1535 -14
rect 1396 -27 1419 -22
rect 1427 -27 1471 -22
rect 1479 -27 1523 -22
rect 1427 -30 1431 -27
rect 1479 -30 1483 -27
rect 1531 -30 1535 -18
rect 1553 -22 1558 44
rect 1572 21 1575 26
rect 1583 17 1587 44
rect 1628 41 1632 44
rect 1660 41 1664 44
rect 1620 14 1624 21
rect 1652 14 1656 21
rect 1610 12 1674 14
rect 1610 8 1612 12
rect 1616 8 1636 12
rect 1640 8 1644 12
rect 1648 8 1668 12
rect 1672 8 1674 12
rect 1610 6 1674 8
rect 1575 -14 1579 -3
rect 1575 -18 1587 -14
rect 1553 -27 1575 -22
rect 1583 -30 1587 -18
rect 1167 -48 1171 -42
rect 1159 -49 1186 -48
rect 1159 -53 1160 -49
rect 1164 -53 1181 -49
rect 1185 -53 1186 -49
rect 1159 -54 1186 -53
rect 1419 -58 1423 -50
rect 1471 -58 1475 -50
rect 1523 -58 1527 -50
rect 1575 -58 1579 -50
rect 1409 -59 1597 -58
rect 1409 -63 1436 -59
rect 1440 -63 1488 -59
rect 1492 -63 1540 -59
rect 1544 -63 1592 -59
rect 1596 -63 1597 -59
rect 1409 -64 1597 -63
rect 1056 -74 1135 -71
rect 1402 -77 1409 -72
rect 1414 -77 1461 -72
rect 1466 -77 1515 -72
rect 1520 -77 1567 -72
rect 446 -145 450 -140
rect 473 -145 477 -140
rect 246 -152 273 -149
rect 246 -156 249 -152
rect 253 -156 266 -152
rect 270 -156 273 -152
rect 246 -158 273 -156
rect 254 -163 258 -158
rect 143 -171 148 -169
rect -19 -176 14 -171
rect 19 -176 148 -171
rect 108 -180 114 -179
rect 108 -184 109 -180
rect 113 -184 114 -180
rect 108 -187 114 -184
rect 143 -187 148 -176
rect 203 -182 212 -179
rect 203 -186 205 -182
rect 209 -186 212 -182
rect 226 -186 239 -183
rect 203 -187 212 -186
rect 108 -191 120 -187
rect 108 -201 114 -191
rect 198 -191 212 -187
rect 140 -199 158 -195
rect 203 -199 212 -191
rect 108 -205 109 -201
rect 113 -205 114 -201
rect 108 -206 114 -205
rect 143 -209 148 -199
rect 203 -203 205 -199
rect 209 -203 212 -199
rect 203 -206 212 -203
rect 218 -209 222 -206
rect 172 -213 222 -209
rect 172 -218 176 -213
rect -24 -223 176 -218
rect 226 -219 230 -206
rect 233 -213 239 -186
rect 262 -213 266 -203
rect 454 -205 458 -185
rect 481 -205 485 -185
rect 728 -148 816 -143
rect 500 -204 527 -201
rect 454 -209 495 -205
rect 429 -211 446 -210
rect 410 -213 446 -211
rect 233 -218 254 -213
rect 262 -218 308 -213
rect 313 -215 446 -213
rect 313 -217 437 -215
rect 313 -218 418 -217
rect -215 -237 -151 -234
rect -215 -241 -212 -237
rect -208 -241 -190 -237
rect -186 -241 -180 -237
rect -176 -241 -158 -237
rect -154 -241 -151 -237
rect -416 -245 -228 -242
rect -215 -243 -151 -241
rect -416 -249 -413 -245
rect -409 -249 -391 -245
rect -387 -249 -361 -245
rect -357 -249 -339 -245
rect -335 -249 -309 -245
rect -305 -249 -287 -245
rect -283 -249 -257 -245
rect -253 -249 -235 -245
rect -231 -249 -228 -245
rect -416 -251 -228 -249
rect -205 -249 -201 -243
rect -173 -249 -169 -243
rect -406 -257 -402 -251
rect -354 -257 -350 -251
rect -302 -257 -298 -251
rect -250 -257 -246 -251
rect -429 -306 -406 -301
rect -429 -372 -424 -306
rect -398 -310 -394 -297
rect -406 -314 -394 -310
rect -376 -306 -354 -301
rect -406 -319 -402 -314
rect -411 -368 -406 -363
rect -398 -372 -394 -359
rect -376 -372 -371 -306
rect -346 -310 -342 -297
rect -294 -301 -290 -297
rect -242 -301 -238 -297
rect -197 -301 -193 -289
rect -165 -301 -161 -289
rect -24 -301 -17 -223
rect -354 -314 -342 -310
rect -324 -306 -302 -301
rect -294 -306 -250 -301
rect -242 -306 -205 -301
rect -197 -306 -173 -301
rect -165 -306 -16 -301
rect -354 -319 -350 -314
rect -359 -368 -354 -363
rect -346 -372 -342 -359
rect -324 -372 -319 -306
rect -305 -329 -302 -324
rect -294 -333 -290 -306
rect -302 -364 -298 -353
rect -302 -368 -290 -364
rect -429 -377 -406 -372
rect -398 -377 -354 -372
rect -346 -377 -302 -372
rect -398 -380 -394 -377
rect -346 -380 -342 -377
rect -294 -380 -290 -368
rect -272 -372 -267 -306
rect -253 -329 -250 -324
rect -242 -333 -238 -306
rect -197 -309 -193 -306
rect -165 -309 -161 -306
rect -154 -307 -16 -306
rect -205 -336 -201 -329
rect -173 -336 -169 -329
rect -215 -338 -151 -336
rect -215 -342 -213 -338
rect -209 -342 -189 -338
rect -185 -342 -181 -338
rect -177 -342 -157 -338
rect -153 -342 -151 -338
rect -215 -344 -151 -342
rect -250 -364 -246 -353
rect -250 -368 -238 -364
rect -272 -377 -250 -372
rect -242 -380 -238 -368
rect -406 -408 -402 -400
rect -354 -408 -350 -400
rect -302 -408 -298 -400
rect -250 -408 -246 -400
rect -416 -409 -228 -408
rect -416 -413 -389 -409
rect -385 -413 -337 -409
rect -333 -413 -285 -409
rect -281 -413 -233 -409
rect -229 -413 -228 -409
rect -416 -414 -228 -413
rect -423 -427 -416 -422
rect -411 -427 -364 -422
rect -359 -427 -310 -422
rect -305 -427 -258 -422
rect 69 -438 74 -223
rect 108 -231 114 -230
rect 108 -235 109 -231
rect 113 -235 114 -231
rect 108 -238 114 -235
rect 143 -238 148 -223
rect 203 -233 212 -230
rect 203 -237 205 -233
rect 209 -237 212 -233
rect 203 -238 212 -237
rect 108 -242 120 -238
rect 108 -252 114 -242
rect 198 -242 212 -238
rect 140 -250 158 -246
rect 203 -250 212 -242
rect 108 -256 109 -252
rect 113 -256 114 -252
rect 108 -257 114 -256
rect 143 -270 148 -250
rect 203 -254 205 -250
rect 209 -254 212 -250
rect 203 -257 212 -254
rect 262 -221 266 -218
rect 473 -219 477 -209
rect 218 -270 222 -239
rect 254 -247 258 -241
rect 246 -248 273 -247
rect 246 -252 247 -248
rect 251 -252 268 -248
rect 272 -252 273 -248
rect 246 -253 273 -252
rect 465 -265 469 -259
rect 490 -265 495 -209
rect 500 -208 503 -204
rect 507 -208 520 -204
rect 524 -208 527 -204
rect 500 -210 527 -208
rect 508 -215 512 -210
rect 516 -265 520 -255
rect 728 -265 733 -148
rect 824 -152 828 -140
rect 816 -156 828 -152
rect 816 -160 820 -156
rect 1625 -163 1689 -160
rect 1625 -167 1628 -163
rect 1632 -167 1650 -163
rect 1654 -167 1660 -163
rect 1664 -167 1682 -163
rect 1686 -167 1689 -163
rect 1154 -173 1181 -170
rect 1154 -177 1157 -173
rect 1161 -177 1174 -173
rect 1178 -177 1181 -173
rect 1424 -171 1612 -168
rect 1625 -169 1689 -167
rect 1424 -175 1427 -171
rect 1431 -175 1449 -171
rect 1453 -175 1479 -171
rect 1483 -175 1501 -171
rect 1505 -175 1531 -171
rect 1535 -175 1553 -171
rect 1557 -175 1583 -171
rect 1587 -175 1605 -171
rect 1609 -175 1612 -171
rect 1424 -177 1612 -175
rect 1635 -175 1639 -169
rect 1667 -175 1671 -169
rect 1154 -179 1181 -177
rect 857 -186 884 -183
rect 1162 -184 1166 -179
rect 1434 -183 1438 -177
rect 1486 -183 1490 -177
rect 1538 -183 1542 -177
rect 1590 -183 1594 -177
rect 857 -190 860 -186
rect 864 -190 877 -186
rect 881 -190 884 -186
rect 857 -192 884 -190
rect 1051 -192 1056 -190
rect 865 -197 869 -192
rect 979 -197 1056 -192
rect 465 -269 479 -265
rect 143 -273 222 -270
rect 473 -270 479 -269
rect 490 -270 508 -265
rect 516 -270 733 -265
rect 757 -251 801 -246
rect 824 -247 828 -240
rect 873 -247 877 -237
rect 429 -278 465 -276
rect 416 -279 465 -278
rect 304 -281 465 -279
rect 304 -284 443 -281
rect 473 -284 477 -270
rect 516 -273 520 -270
rect 163 -296 217 -293
rect 163 -300 166 -296
rect 170 -300 183 -296
rect 187 -300 193 -296
rect 197 -300 210 -296
rect 214 -300 217 -296
rect 163 -302 217 -300
rect 171 -307 175 -302
rect 198 -307 202 -302
rect 508 -299 512 -293
rect 500 -300 527 -299
rect 500 -304 501 -300
rect 505 -304 522 -300
rect 526 -304 527 -300
rect 500 -305 527 -304
rect 465 -330 469 -324
rect 457 -331 484 -330
rect 457 -335 458 -331
rect 462 -335 479 -331
rect 483 -335 484 -331
rect 457 -336 484 -335
rect 179 -367 183 -347
rect 206 -367 210 -347
rect 225 -366 252 -363
rect 179 -371 220 -367
rect 107 -377 171 -372
rect 198 -381 202 -371
rect 190 -427 194 -421
rect 215 -427 220 -371
rect 225 -370 228 -366
rect 232 -370 245 -366
rect 249 -370 252 -366
rect 225 -372 252 -370
rect 233 -377 237 -372
rect 241 -427 245 -417
rect 757 -424 762 -251
rect 824 -252 865 -247
rect 873 -252 936 -247
rect 979 -252 984 -197
rect 1016 -201 1022 -200
rect 1016 -205 1017 -201
rect 1021 -205 1022 -201
rect 1016 -208 1022 -205
rect 1051 -208 1056 -197
rect 1111 -203 1120 -200
rect 1111 -207 1113 -203
rect 1117 -207 1120 -203
rect 1134 -207 1147 -204
rect 1111 -208 1120 -207
rect 1016 -212 1028 -208
rect 1016 -222 1022 -212
rect 1106 -212 1120 -208
rect 1048 -220 1066 -216
rect 1111 -220 1120 -212
rect 1016 -226 1017 -222
rect 1021 -226 1022 -222
rect 1016 -227 1022 -226
rect 1051 -230 1056 -220
rect 1111 -224 1113 -220
rect 1117 -224 1120 -220
rect 1111 -227 1120 -224
rect 1126 -230 1130 -227
rect 1080 -234 1130 -230
rect 1080 -239 1084 -234
rect 824 -255 828 -252
rect 873 -255 877 -252
rect 809 -259 846 -255
rect 809 -265 813 -259
rect 842 -265 846 -259
rect 926 -257 984 -252
rect 993 -244 1084 -239
rect 1134 -240 1138 -227
rect 1141 -234 1147 -207
rect 1170 -234 1174 -224
rect 1411 -232 1434 -227
rect 1220 -234 1229 -233
rect 1141 -239 1162 -234
rect 1170 -239 1229 -234
rect 865 -281 869 -275
rect 857 -282 884 -281
rect 801 -291 805 -285
rect 834 -291 838 -285
rect 857 -286 858 -282
rect 862 -286 879 -282
rect 883 -286 884 -282
rect 857 -287 884 -286
rect 793 -292 820 -291
rect 793 -296 794 -292
rect 798 -296 815 -292
rect 819 -296 820 -292
rect 793 -297 820 -296
rect 826 -292 853 -291
rect 826 -296 827 -292
rect 831 -296 848 -292
rect 852 -296 853 -292
rect 826 -297 853 -296
rect 429 -427 762 -424
rect 190 -431 204 -427
rect 198 -432 204 -431
rect 215 -432 233 -427
rect 241 -432 317 -427
rect 322 -429 762 -427
rect 322 -432 440 -429
rect 69 -443 190 -438
rect 198 -446 202 -432
rect 241 -435 245 -432
rect 413 -433 440 -432
rect 429 -455 936 -453
rect 233 -461 237 -455
rect 415 -456 936 -455
rect 331 -458 936 -456
rect 993 -458 998 -244
rect 1016 -252 1022 -251
rect 1016 -256 1017 -252
rect 1021 -256 1022 -252
rect 1016 -259 1022 -256
rect 1051 -259 1056 -244
rect 1111 -254 1120 -251
rect 1111 -258 1113 -254
rect 1117 -258 1120 -254
rect 1111 -259 1120 -258
rect 1016 -263 1028 -259
rect 1016 -273 1022 -263
rect 1106 -263 1120 -259
rect 1048 -271 1066 -267
rect 1111 -271 1120 -263
rect 1016 -277 1017 -273
rect 1021 -277 1022 -273
rect 1016 -278 1022 -277
rect 1051 -291 1056 -271
rect 1111 -275 1113 -271
rect 1117 -275 1120 -271
rect 1111 -278 1120 -275
rect 1170 -242 1174 -239
rect 1126 -291 1130 -260
rect 1162 -268 1166 -262
rect 1154 -269 1181 -268
rect 1154 -273 1155 -269
rect 1159 -273 1176 -269
rect 1180 -273 1181 -269
rect 1154 -274 1181 -273
rect 1220 -278 1229 -239
rect 1411 -278 1416 -232
rect 1442 -236 1446 -223
rect 1220 -283 1416 -278
rect 1220 -284 1229 -283
rect 1051 -294 1130 -291
rect 1411 -298 1416 -283
rect 1434 -240 1446 -236
rect 1464 -232 1486 -227
rect 1434 -245 1438 -240
rect 1429 -294 1434 -289
rect 1442 -298 1446 -285
rect 1464 -298 1469 -232
rect 1494 -236 1498 -223
rect 1546 -227 1550 -223
rect 1598 -227 1602 -223
rect 1643 -227 1647 -215
rect 1675 -227 1679 -215
rect 1486 -240 1498 -236
rect 1516 -232 1538 -227
rect 1546 -232 1590 -227
rect 1598 -232 1635 -227
rect 1643 -232 1667 -227
rect 1675 -232 1689 -227
rect 1486 -245 1490 -240
rect 1481 -294 1486 -289
rect 1494 -298 1498 -285
rect 1516 -298 1521 -232
rect 1535 -255 1538 -250
rect 1546 -259 1550 -232
rect 1538 -290 1542 -279
rect 1538 -294 1550 -290
rect 1411 -303 1434 -298
rect 1442 -303 1486 -298
rect 1494 -303 1538 -298
rect 1442 -306 1446 -303
rect 1494 -306 1498 -303
rect 1546 -306 1550 -294
rect 1568 -298 1573 -232
rect 1587 -255 1590 -250
rect 1598 -259 1602 -232
rect 1643 -235 1647 -232
rect 1675 -235 1679 -232
rect 1635 -262 1639 -255
rect 1667 -262 1671 -255
rect 1625 -264 1689 -262
rect 1625 -268 1627 -264
rect 1631 -268 1651 -264
rect 1655 -268 1659 -264
rect 1663 -268 1683 -264
rect 1687 -268 1689 -264
rect 1625 -270 1689 -268
rect 1590 -290 1594 -279
rect 1590 -294 1602 -290
rect 1568 -303 1590 -298
rect 1598 -306 1602 -294
rect 1434 -334 1438 -326
rect 1486 -334 1490 -326
rect 1538 -334 1542 -326
rect 1590 -334 1594 -326
rect 1424 -335 1612 -334
rect 1424 -339 1451 -335
rect 1455 -339 1503 -335
rect 1507 -339 1555 -335
rect 1559 -339 1607 -335
rect 1611 -339 1612 -335
rect 1424 -340 1612 -339
rect 1417 -353 1424 -348
rect 1429 -353 1476 -348
rect 1481 -353 1530 -348
rect 1535 -353 1582 -348
rect 331 -461 442 -458
rect 225 -462 252 -461
rect 225 -466 226 -462
rect 230 -466 247 -462
rect 251 -466 252 -462
rect 926 -463 998 -458
rect 225 -467 252 -466
rect 190 -492 194 -486
rect 182 -493 209 -492
rect 182 -497 183 -493
rect 187 -497 204 -493
rect 208 -497 209 -493
rect 182 -498 209 -497
rect 952 -696 979 -693
rect 952 -700 955 -696
rect 959 -700 972 -696
rect 976 -700 979 -696
rect 952 -702 979 -700
rect 1203 -698 1230 -695
rect 1203 -702 1206 -698
rect 1210 -702 1223 -698
rect 1227 -702 1230 -698
rect 960 -707 964 -702
rect 1203 -704 1230 -702
rect 423 -735 891 -730
rect 423 -752 431 -735
rect 335 -757 433 -752
rect -118 -819 -54 -816
rect -118 -823 -115 -819
rect -111 -823 -93 -819
rect -89 -823 -83 -819
rect -79 -823 -61 -819
rect -57 -823 -54 -819
rect -319 -827 -131 -824
rect -118 -825 -54 -823
rect -319 -831 -316 -827
rect -312 -831 -294 -827
rect -290 -831 -264 -827
rect -260 -831 -242 -827
rect -238 -831 -212 -827
rect -208 -831 -190 -827
rect -186 -831 -160 -827
rect -156 -831 -138 -827
rect -134 -831 -131 -827
rect -319 -833 -131 -831
rect -108 -831 -104 -825
rect -76 -831 -72 -825
rect -309 -839 -305 -833
rect -257 -839 -253 -833
rect -205 -839 -201 -833
rect -153 -839 -149 -833
rect 335 -859 340 -757
rect 375 -759 433 -757
rect 423 -761 431 -759
rect 618 -785 672 -782
rect 618 -789 621 -785
rect 625 -789 638 -785
rect 642 -789 648 -785
rect 652 -789 665 -785
rect 669 -789 672 -785
rect 618 -791 672 -789
rect 879 -789 891 -735
rect 879 -790 929 -789
rect 626 -796 630 -791
rect 653 -796 657 -791
rect 879 -795 960 -790
rect 968 -799 972 -787
rect 1211 -709 1215 -704
rect 634 -856 638 -836
rect 661 -856 665 -836
rect 960 -803 972 -799
rect 1132 -797 1211 -792
rect 960 -807 964 -803
rect 680 -855 707 -852
rect 634 -860 675 -856
rect 335 -867 340 -864
rect 423 -866 626 -861
rect -332 -888 -309 -883
rect -332 -954 -327 -888
rect -301 -892 -297 -879
rect -309 -896 -297 -892
rect -279 -888 -257 -883
rect -309 -901 -305 -896
rect -314 -950 -309 -945
rect -301 -954 -297 -941
rect -279 -954 -274 -888
rect -249 -892 -245 -879
rect -197 -883 -193 -879
rect -145 -883 -141 -879
rect -100 -883 -96 -871
rect -68 -883 -64 -871
rect -257 -896 -245 -892
rect -227 -888 -205 -883
rect -197 -888 -153 -883
rect -145 -888 -108 -883
rect -100 -888 -76 -883
rect -68 -884 -7 -883
rect -68 -888 -6 -884
rect 322 -884 382 -883
rect 424 -884 429 -866
rect 653 -870 657 -860
rect 322 -888 429 -884
rect -257 -901 -253 -896
rect -262 -950 -257 -945
rect -249 -954 -245 -941
rect -227 -954 -222 -888
rect -208 -911 -205 -906
rect -197 -915 -193 -888
rect -205 -946 -201 -935
rect -205 -950 -193 -946
rect -332 -959 -309 -954
rect -301 -959 -257 -954
rect -249 -959 -205 -954
rect -301 -962 -297 -959
rect -249 -962 -245 -959
rect -197 -962 -193 -950
rect -175 -954 -170 -888
rect -156 -911 -153 -906
rect -145 -915 -141 -888
rect -100 -891 -96 -888
rect -68 -891 -64 -888
rect -57 -890 -6 -888
rect -108 -918 -104 -911
rect -76 -918 -72 -911
rect -118 -920 -54 -918
rect -118 -924 -116 -920
rect -112 -924 -92 -920
rect -88 -924 -84 -920
rect -80 -924 -60 -920
rect -56 -924 -54 -920
rect -118 -926 -54 -924
rect -153 -946 -149 -935
rect -153 -950 -141 -946
rect -175 -959 -153 -954
rect -145 -962 -141 -950
rect -14 -957 -6 -890
rect 645 -916 649 -910
rect 670 -916 675 -860
rect 680 -859 683 -855
rect 687 -859 700 -855
rect 704 -859 707 -855
rect 680 -861 707 -859
rect 688 -866 692 -861
rect 1001 -833 1028 -830
rect 1001 -837 1004 -833
rect 1008 -837 1021 -833
rect 1025 -837 1028 -833
rect 1001 -839 1028 -837
rect 1009 -844 1013 -839
rect 696 -916 700 -906
rect 874 -893 938 -887
rect 874 -898 945 -893
rect 968 -894 972 -887
rect 1017 -894 1021 -884
rect 1132 -894 1137 -797
rect 1219 -801 1223 -789
rect 1211 -805 1223 -801
rect 1211 -809 1215 -805
rect 1252 -835 1279 -832
rect 1252 -839 1255 -835
rect 1259 -839 1272 -835
rect 1276 -839 1279 -835
rect 1252 -841 1279 -839
rect 2009 -836 2073 -833
rect 2009 -840 2012 -836
rect 2016 -840 2034 -836
rect 2038 -840 2044 -836
rect 2048 -840 2066 -836
rect 2070 -840 2073 -836
rect 1260 -846 1264 -841
rect 1808 -844 1996 -841
rect 2009 -842 2073 -840
rect 1808 -848 1811 -844
rect 1815 -848 1833 -844
rect 1837 -848 1863 -844
rect 1867 -848 1885 -844
rect 1889 -848 1915 -844
rect 1919 -848 1937 -844
rect 1941 -848 1967 -844
rect 1971 -848 1989 -844
rect 1993 -848 1996 -844
rect 1808 -850 1996 -848
rect 2019 -848 2023 -842
rect 2051 -848 2055 -842
rect 874 -916 882 -898
rect 968 -899 1009 -894
rect 1017 -899 1137 -894
rect 968 -902 972 -899
rect 1017 -902 1021 -899
rect 953 -906 990 -902
rect 953 -912 957 -906
rect 986 -912 990 -906
rect 645 -920 659 -916
rect 653 -921 659 -920
rect 670 -921 688 -916
rect 696 -921 882 -916
rect 580 -932 645 -927
rect 234 -938 261 -935
rect 234 -942 237 -938
rect 241 -942 254 -938
rect 258 -942 261 -938
rect 234 -944 261 -942
rect 242 -949 246 -944
rect 131 -957 136 -955
rect -15 -962 2 -957
rect 7 -962 136 -957
rect 96 -966 102 -965
rect 96 -970 97 -966
rect 101 -970 102 -966
rect 96 -973 102 -970
rect 131 -973 136 -962
rect 191 -968 200 -965
rect 191 -972 193 -968
rect 197 -972 200 -968
rect 214 -972 227 -969
rect 191 -973 200 -972
rect 96 -977 108 -973
rect -309 -990 -305 -982
rect -257 -990 -253 -982
rect -205 -990 -201 -982
rect -153 -990 -149 -982
rect 96 -987 102 -977
rect 186 -977 200 -973
rect 128 -985 146 -981
rect 191 -985 200 -977
rect -319 -991 -131 -990
rect -319 -995 -292 -991
rect -288 -995 -240 -991
rect -236 -995 -188 -991
rect -184 -995 -136 -991
rect -132 -995 -131 -991
rect 96 -991 97 -987
rect 101 -991 102 -987
rect 96 -992 102 -991
rect -319 -996 -131 -995
rect 131 -995 136 -985
rect 191 -989 193 -985
rect 197 -989 200 -985
rect 191 -992 200 -989
rect 206 -995 210 -992
rect 160 -999 210 -995
rect -31 -1004 -25 -1003
rect 160 -1004 164 -999
rect -326 -1009 -319 -1004
rect -314 -1009 -267 -1004
rect -262 -1009 -213 -1004
rect -208 -1009 -161 -1004
rect -31 -1009 164 -1004
rect 214 -1005 218 -992
rect 221 -999 227 -972
rect 580 -977 585 -932
rect 653 -935 657 -921
rect 696 -924 700 -921
rect 874 -924 882 -921
rect 250 -999 254 -989
rect 423 -982 585 -977
rect 1163 -900 1196 -895
rect 1219 -896 1223 -889
rect 1268 -896 1272 -886
rect 1818 -856 1822 -850
rect 1870 -856 1874 -850
rect 1922 -856 1926 -850
rect 1974 -856 1978 -850
rect 1009 -928 1013 -922
rect 1001 -929 1028 -928
rect 945 -938 949 -932
rect 978 -938 982 -932
rect 1001 -933 1002 -929
rect 1006 -933 1023 -929
rect 1027 -933 1028 -929
rect 1001 -934 1028 -933
rect 937 -939 964 -938
rect 937 -943 938 -939
rect 942 -943 959 -939
rect 963 -943 964 -939
rect 937 -944 964 -943
rect 970 -939 997 -938
rect 970 -943 971 -939
rect 975 -943 992 -939
rect 996 -943 997 -939
rect 970 -944 997 -943
rect 688 -950 692 -944
rect 680 -951 707 -950
rect 680 -955 681 -951
rect 685 -955 702 -951
rect 706 -955 707 -951
rect 680 -956 707 -955
rect 645 -981 649 -975
rect 637 -982 664 -981
rect 423 -999 428 -982
rect 637 -986 638 -982
rect 642 -986 659 -982
rect 663 -986 664 -982
rect 637 -987 664 -986
rect 221 -1004 242 -999
rect 250 -1004 326 -999
rect 331 -1004 428 -999
rect -137 -1042 -73 -1039
rect -137 -1046 -134 -1042
rect -130 -1046 -112 -1042
rect -108 -1046 -102 -1042
rect -98 -1046 -80 -1042
rect -76 -1046 -73 -1042
rect -338 -1050 -150 -1047
rect -137 -1048 -73 -1046
rect -338 -1054 -335 -1050
rect -331 -1054 -313 -1050
rect -309 -1054 -283 -1050
rect -279 -1054 -261 -1050
rect -257 -1054 -231 -1050
rect -227 -1054 -209 -1050
rect -205 -1054 -179 -1050
rect -175 -1054 -157 -1050
rect -153 -1054 -150 -1050
rect -338 -1056 -150 -1054
rect -127 -1054 -123 -1048
rect -95 -1054 -91 -1048
rect -328 -1062 -324 -1056
rect -276 -1062 -272 -1056
rect -224 -1062 -220 -1056
rect -172 -1062 -168 -1056
rect -351 -1111 -328 -1106
rect -3297 -1145 -3270 -1142
rect -3297 -1149 -3294 -1145
rect -3290 -1149 -3277 -1145
rect -3273 -1149 -3270 -1145
rect -3297 -1151 -3270 -1149
rect -3289 -1156 -3285 -1151
rect -3453 -1172 -3426 -1169
rect -3453 -1176 -3450 -1172
rect -3446 -1176 -3433 -1172
rect -3429 -1176 -3426 -1172
rect -3453 -1178 -3426 -1176
rect -3445 -1183 -3441 -1178
rect -3556 -1191 -3551 -1189
rect -3591 -1196 -3551 -1191
rect -3591 -1200 -3585 -1199
rect -3591 -1204 -3590 -1200
rect -3586 -1204 -3585 -1200
rect -3591 -1207 -3585 -1204
rect -3556 -1207 -3551 -1196
rect -3496 -1202 -3487 -1199
rect -3496 -1206 -3494 -1202
rect -3490 -1206 -3487 -1202
rect -3473 -1206 -3460 -1203
rect -3496 -1207 -3487 -1206
rect -3591 -1211 -3579 -1207
rect -3591 -1221 -3585 -1211
rect -3501 -1211 -3487 -1207
rect -3559 -1219 -3541 -1215
rect -3496 -1219 -3487 -1211
rect -3591 -1225 -3590 -1221
rect -3586 -1225 -3585 -1221
rect -3591 -1226 -3585 -1225
rect -3556 -1229 -3551 -1219
rect -3496 -1223 -3494 -1219
rect -3490 -1223 -3487 -1219
rect -3496 -1226 -3487 -1223
rect -3481 -1229 -3477 -1226
rect -3527 -1233 -3477 -1229
rect -3527 -1238 -3523 -1233
rect -3591 -1243 -3523 -1238
rect -3473 -1239 -3469 -1226
rect -3466 -1233 -3460 -1206
rect -3362 -1188 -3335 -1185
rect -3362 -1192 -3359 -1188
rect -3355 -1192 -3342 -1188
rect -3338 -1192 -3335 -1188
rect -3362 -1194 -3335 -1192
rect -3437 -1233 -3433 -1223
rect -3354 -1199 -3350 -1194
rect -3466 -1238 -3445 -1233
rect -3437 -1238 -3426 -1233
rect -3591 -1251 -3585 -1250
rect -3591 -1255 -3590 -1251
rect -3586 -1255 -3585 -1251
rect -3591 -1258 -3585 -1255
rect -3556 -1258 -3551 -1243
rect -3496 -1253 -3487 -1250
rect -3496 -1257 -3494 -1253
rect -3490 -1257 -3487 -1253
rect -3496 -1258 -3487 -1257
rect -3591 -1262 -3579 -1258
rect -3591 -1272 -3585 -1262
rect -3501 -1262 -3487 -1258
rect -3559 -1270 -3541 -1266
rect -3496 -1270 -3487 -1262
rect -3591 -1276 -3590 -1272
rect -3586 -1276 -3585 -1272
rect -3591 -1277 -3585 -1276
rect -3556 -1290 -3551 -1270
rect -3496 -1274 -3494 -1270
rect -3490 -1274 -3487 -1270
rect -3496 -1277 -3487 -1274
rect -3437 -1241 -3433 -1238
rect -3188 -1157 -3134 -1154
rect -3188 -1161 -3185 -1157
rect -3181 -1161 -3168 -1157
rect -3164 -1161 -3158 -1157
rect -3154 -1161 -3141 -1157
rect -3137 -1161 -3134 -1157
rect -3188 -1163 -3134 -1161
rect -3180 -1168 -3176 -1163
rect -3153 -1168 -3149 -1163
rect -351 -1177 -346 -1111
rect -320 -1115 -316 -1102
rect -328 -1119 -316 -1115
rect -298 -1111 -276 -1106
rect -328 -1124 -324 -1119
rect -333 -1173 -328 -1168
rect -320 -1177 -316 -1164
rect -298 -1177 -293 -1111
rect -268 -1115 -264 -1102
rect -216 -1106 -212 -1102
rect -164 -1106 -160 -1102
rect -119 -1106 -115 -1094
rect -87 -1106 -83 -1094
rect -31 -1106 -25 -1009
rect -276 -1119 -264 -1115
rect -246 -1111 -224 -1106
rect -216 -1111 -172 -1106
rect -164 -1111 -127 -1106
rect -119 -1111 -95 -1106
rect -87 -1111 -23 -1106
rect -276 -1124 -272 -1119
rect -281 -1173 -276 -1168
rect -268 -1177 -264 -1164
rect -246 -1177 -241 -1111
rect -227 -1134 -224 -1129
rect -216 -1138 -212 -1111
rect -224 -1169 -220 -1158
rect -224 -1173 -212 -1169
rect -351 -1182 -328 -1177
rect -320 -1182 -276 -1177
rect -268 -1182 -224 -1177
rect -320 -1185 -316 -1182
rect -268 -1185 -264 -1182
rect -216 -1185 -212 -1173
rect -194 -1177 -189 -1111
rect -175 -1134 -172 -1129
rect -164 -1138 -160 -1111
rect -119 -1114 -115 -1111
rect -87 -1114 -83 -1111
rect -77 -1112 -23 -1111
rect -127 -1141 -123 -1134
rect -95 -1141 -91 -1134
rect -137 -1143 -73 -1141
rect -137 -1147 -135 -1143
rect -131 -1147 -111 -1143
rect -107 -1147 -103 -1143
rect -99 -1147 -79 -1143
rect -75 -1147 -73 -1143
rect -137 -1149 -73 -1147
rect -172 -1169 -168 -1158
rect -172 -1173 -160 -1169
rect -194 -1182 -172 -1177
rect -164 -1185 -160 -1173
rect -3172 -1228 -3168 -1208
rect -3145 -1228 -3141 -1208
rect -328 -1213 -324 -1205
rect -276 -1213 -272 -1205
rect -224 -1213 -220 -1205
rect -172 -1213 -168 -1205
rect -338 -1214 -150 -1213
rect -338 -1218 -311 -1214
rect -307 -1218 -259 -1214
rect -255 -1218 -207 -1214
rect -203 -1218 -155 -1214
rect -151 -1218 -150 -1214
rect -338 -1219 -150 -1218
rect 57 -1224 62 -1009
rect 96 -1017 102 -1016
rect 96 -1021 97 -1017
rect 101 -1021 102 -1017
rect 96 -1024 102 -1021
rect 131 -1024 136 -1009
rect 191 -1019 200 -1016
rect 191 -1023 193 -1019
rect 197 -1023 200 -1019
rect 191 -1024 200 -1023
rect 96 -1028 108 -1024
rect 96 -1038 102 -1028
rect 186 -1028 200 -1024
rect 128 -1036 146 -1032
rect 191 -1036 200 -1028
rect 96 -1042 97 -1038
rect 101 -1042 102 -1038
rect 96 -1043 102 -1042
rect 131 -1056 136 -1036
rect 191 -1040 193 -1036
rect 197 -1040 200 -1036
rect 191 -1043 200 -1040
rect 250 -1007 254 -1004
rect 375 -1005 428 -1004
rect 206 -1056 210 -1025
rect 242 -1033 246 -1027
rect 541 -1030 595 -1027
rect 234 -1034 261 -1033
rect 234 -1038 235 -1034
rect 239 -1038 256 -1034
rect 260 -1038 261 -1034
rect 541 -1034 544 -1030
rect 548 -1034 561 -1030
rect 565 -1034 571 -1030
rect 575 -1034 588 -1030
rect 592 -1034 595 -1030
rect 541 -1036 595 -1034
rect 759 -1030 813 -1027
rect 759 -1034 762 -1030
rect 766 -1034 779 -1030
rect 783 -1034 789 -1030
rect 793 -1034 806 -1030
rect 810 -1034 813 -1030
rect 759 -1036 813 -1034
rect 234 -1039 261 -1038
rect 131 -1059 210 -1056
rect 549 -1041 553 -1036
rect 576 -1041 580 -1036
rect 767 -1041 771 -1036
rect 794 -1041 798 -1036
rect 151 -1082 205 -1079
rect 151 -1086 154 -1082
rect 158 -1086 171 -1082
rect 175 -1086 181 -1082
rect 185 -1086 198 -1082
rect 202 -1086 205 -1082
rect 151 -1088 205 -1086
rect 159 -1093 163 -1088
rect 186 -1093 190 -1088
rect 557 -1101 561 -1081
rect 584 -1101 588 -1081
rect 603 -1100 630 -1097
rect 404 -1106 413 -1104
rect 557 -1105 598 -1101
rect 404 -1111 549 -1106
rect 404 -1128 413 -1111
rect 576 -1115 580 -1105
rect 423 -1119 537 -1118
rect 304 -1129 413 -1128
rect 422 -1123 537 -1119
rect 304 -1133 414 -1129
rect 167 -1153 171 -1133
rect 194 -1153 198 -1133
rect 422 -1140 428 -1123
rect 313 -1145 428 -1140
rect 213 -1152 240 -1149
rect 167 -1157 208 -1153
rect 95 -1163 159 -1158
rect 186 -1167 190 -1157
rect 178 -1213 182 -1207
rect 203 -1213 208 -1157
rect 213 -1156 216 -1152
rect 220 -1156 233 -1152
rect 237 -1156 240 -1152
rect 213 -1158 240 -1156
rect 221 -1163 225 -1158
rect 532 -1172 537 -1123
rect 568 -1161 572 -1155
rect 593 -1161 598 -1105
rect 603 -1104 606 -1100
rect 610 -1104 623 -1100
rect 627 -1104 630 -1100
rect 603 -1106 630 -1104
rect 775 -1101 779 -1081
rect 802 -1101 806 -1081
rect 821 -1100 848 -1097
rect 775 -1105 816 -1101
rect 723 -1106 755 -1105
rect 611 -1111 615 -1106
rect 663 -1111 767 -1106
rect 619 -1161 623 -1151
rect 663 -1161 668 -1111
rect 794 -1115 798 -1105
rect 568 -1165 582 -1161
rect 576 -1166 582 -1165
rect 593 -1166 611 -1161
rect 619 -1166 668 -1161
rect 786 -1161 790 -1155
rect 811 -1161 816 -1105
rect 821 -1104 824 -1100
rect 828 -1104 841 -1100
rect 845 -1104 848 -1100
rect 821 -1106 848 -1104
rect 868 -1105 934 -1102
rect 1163 -1105 1168 -900
rect 1219 -901 1260 -896
rect 1268 -901 1376 -896
rect 1219 -904 1223 -901
rect 1268 -904 1272 -901
rect 1204 -908 1241 -904
rect 1204 -914 1208 -908
rect 1237 -914 1241 -908
rect 1371 -922 1376 -901
rect 1606 -903 1633 -900
rect 1606 -907 1609 -903
rect 1613 -907 1626 -903
rect 1630 -907 1633 -903
rect 1606 -909 1633 -907
rect 1795 -905 1818 -900
rect 1614 -914 1618 -909
rect 1503 -922 1508 -920
rect 1260 -930 1264 -924
rect 1371 -927 1508 -922
rect 1252 -931 1279 -930
rect 1196 -940 1200 -934
rect 1229 -940 1233 -934
rect 1252 -935 1253 -931
rect 1257 -935 1274 -931
rect 1278 -935 1279 -931
rect 1252 -936 1279 -935
rect 1468 -931 1474 -930
rect 1468 -935 1469 -931
rect 1473 -935 1474 -931
rect 1468 -938 1474 -935
rect 1503 -938 1508 -927
rect 1563 -933 1572 -930
rect 1563 -937 1565 -933
rect 1569 -937 1572 -933
rect 1586 -937 1599 -934
rect 1563 -938 1572 -937
rect 1188 -941 1215 -940
rect 1188 -945 1189 -941
rect 1193 -945 1210 -941
rect 1214 -945 1215 -941
rect 1188 -946 1215 -945
rect 1221 -941 1248 -940
rect 1221 -945 1222 -941
rect 1226 -945 1243 -941
rect 1247 -945 1248 -941
rect 1221 -946 1248 -945
rect 1468 -942 1480 -938
rect 1468 -952 1474 -942
rect 1558 -942 1572 -938
rect 1500 -950 1518 -946
rect 1563 -950 1572 -942
rect 1468 -956 1469 -952
rect 1473 -956 1474 -952
rect 1468 -957 1474 -956
rect 1503 -960 1508 -950
rect 1563 -954 1565 -950
rect 1569 -954 1572 -950
rect 1563 -957 1572 -954
rect 1578 -960 1582 -957
rect 1532 -964 1582 -960
rect 829 -1111 833 -1106
rect 868 -1110 1168 -1105
rect 1245 -969 1251 -968
rect 1532 -969 1536 -964
rect 1245 -974 1536 -969
rect 1586 -970 1590 -957
rect 1593 -964 1599 -937
rect 1795 -937 1800 -905
rect 1826 -909 1830 -896
rect 1622 -964 1626 -954
rect 1765 -942 1800 -937
rect 1765 -964 1771 -942
rect 1593 -969 1614 -964
rect 1622 -969 1771 -964
rect 837 -1161 841 -1151
rect 868 -1113 934 -1110
rect 868 -1161 879 -1113
rect 786 -1165 800 -1161
rect 794 -1166 800 -1165
rect 811 -1166 829 -1161
rect 837 -1166 881 -1161
rect 532 -1177 568 -1172
rect 576 -1180 580 -1166
rect 619 -1169 623 -1166
rect 229 -1213 233 -1203
rect 178 -1217 192 -1213
rect 186 -1218 192 -1217
rect 203 -1218 221 -1213
rect 229 -1218 335 -1213
rect 340 -1218 347 -1213
rect -3126 -1227 -3099 -1224
rect -3172 -1232 -3131 -1228
rect -3481 -1290 -3477 -1259
rect -3346 -1249 -3342 -1239
rect -3306 -1244 -3289 -1239
rect -3281 -1248 -3277 -1236
rect -3187 -1238 -3180 -1233
rect -3153 -1242 -3149 -1232
rect -3362 -1254 -3354 -1249
rect -3346 -1254 -3333 -1249
rect -3289 -1252 -3277 -1248
rect -3346 -1257 -3342 -1254
rect -3445 -1267 -3441 -1261
rect -3453 -1268 -3426 -1267
rect -3453 -1272 -3452 -1268
rect -3448 -1272 -3431 -1268
rect -3427 -1272 -3426 -1268
rect -3453 -1273 -3426 -1272
rect -3289 -1256 -3285 -1252
rect -3354 -1283 -3350 -1277
rect -3362 -1284 -3335 -1283
rect -3362 -1288 -3361 -1284
rect -3357 -1288 -3340 -1284
rect -3336 -1288 -3335 -1284
rect -3362 -1289 -3335 -1288
rect -3556 -1293 -3477 -1290
rect -3248 -1282 -3221 -1279
rect -3248 -1286 -3245 -1282
rect -3241 -1286 -3228 -1282
rect -3224 -1286 -3221 -1282
rect -3248 -1288 -3221 -1286
rect -3161 -1288 -3157 -1282
rect -3136 -1288 -3131 -1232
rect -3126 -1231 -3123 -1227
rect -3119 -1231 -3106 -1227
rect -3102 -1231 -3099 -1227
rect -3126 -1233 -3099 -1231
rect -345 -1232 -338 -1227
rect -333 -1232 -286 -1227
rect -281 -1232 -232 -1227
rect -227 -1232 -180 -1227
rect 57 -1229 178 -1224
rect 186 -1232 190 -1218
rect 229 -1221 233 -1218
rect -3118 -1238 -3114 -1233
rect 679 -1177 786 -1172
rect 611 -1195 615 -1189
rect 603 -1196 630 -1195
rect 603 -1200 604 -1196
rect 608 -1200 625 -1196
rect 629 -1200 630 -1196
rect 603 -1201 630 -1200
rect 568 -1226 572 -1220
rect 560 -1227 587 -1226
rect 560 -1231 561 -1227
rect 565 -1231 582 -1227
rect 586 -1231 587 -1227
rect 560 -1232 587 -1231
rect 221 -1247 225 -1241
rect 679 -1244 684 -1177
rect 794 -1180 798 -1166
rect 837 -1169 841 -1166
rect 868 -1167 879 -1166
rect 829 -1195 833 -1189
rect 821 -1196 848 -1195
rect 821 -1200 822 -1196
rect 826 -1200 843 -1196
rect 847 -1200 848 -1196
rect 821 -1201 848 -1200
rect 871 -1210 929 -1209
rect 1245 -1210 1251 -974
rect 1468 -982 1474 -981
rect 1468 -986 1469 -982
rect 1473 -986 1474 -982
rect 1468 -989 1474 -986
rect 1503 -989 1508 -974
rect 1563 -984 1572 -981
rect 1563 -988 1565 -984
rect 1569 -988 1572 -984
rect 1563 -989 1572 -988
rect 1468 -993 1480 -989
rect 1468 -1003 1474 -993
rect 1558 -993 1572 -989
rect 1500 -1001 1518 -997
rect 1563 -1001 1572 -993
rect 1468 -1007 1469 -1003
rect 1473 -1007 1474 -1003
rect 1468 -1008 1474 -1007
rect 1503 -1021 1508 -1001
rect 1563 -1005 1565 -1001
rect 1569 -1005 1572 -1001
rect 1563 -1008 1572 -1005
rect 1622 -972 1626 -969
rect 1578 -1021 1582 -990
rect 1795 -971 1800 -942
rect 1818 -913 1830 -909
rect 1848 -905 1870 -900
rect 1818 -918 1822 -913
rect 1813 -967 1818 -962
rect 1826 -971 1830 -958
rect 1848 -971 1853 -905
rect 1878 -909 1882 -896
rect 1930 -900 1934 -896
rect 1982 -900 1986 -896
rect 2027 -900 2031 -888
rect 2059 -900 2063 -888
rect 1870 -913 1882 -909
rect 1900 -905 1922 -900
rect 1930 -905 1974 -900
rect 1982 -905 2019 -900
rect 2027 -905 2051 -900
rect 2059 -905 2073 -900
rect 1870 -918 1874 -913
rect 1865 -967 1870 -962
rect 1878 -971 1882 -958
rect 1900 -971 1905 -905
rect 1919 -928 1922 -923
rect 1930 -932 1934 -905
rect 1922 -963 1926 -952
rect 1922 -967 1934 -963
rect 1795 -976 1818 -971
rect 1826 -976 1870 -971
rect 1878 -976 1922 -971
rect 1826 -979 1830 -976
rect 1878 -979 1882 -976
rect 1930 -979 1934 -967
rect 1952 -971 1957 -905
rect 1971 -928 1974 -923
rect 1982 -932 1986 -905
rect 2027 -908 2031 -905
rect 2059 -908 2063 -905
rect 2019 -935 2023 -928
rect 2051 -935 2055 -928
rect 2009 -937 2073 -935
rect 2009 -941 2011 -937
rect 2015 -941 2035 -937
rect 2039 -941 2043 -937
rect 2047 -941 2067 -937
rect 2071 -941 2073 -937
rect 2009 -943 2073 -941
rect 1974 -963 1978 -952
rect 1974 -967 1986 -963
rect 1952 -976 1974 -971
rect 1982 -979 1986 -967
rect 1614 -998 1618 -992
rect 1606 -999 1633 -998
rect 1606 -1003 1607 -999
rect 1611 -1003 1628 -999
rect 1632 -1003 1633 -999
rect 1606 -1004 1633 -1003
rect 1818 -1007 1822 -999
rect 1870 -1007 1874 -999
rect 1922 -1007 1926 -999
rect 1974 -1007 1978 -999
rect 1808 -1008 1996 -1007
rect 1808 -1012 1835 -1008
rect 1839 -1012 1887 -1008
rect 1891 -1012 1939 -1008
rect 1943 -1012 1991 -1008
rect 1995 -1012 1996 -1008
rect 1808 -1013 1996 -1012
rect 1503 -1024 1582 -1021
rect 1801 -1026 1808 -1021
rect 1813 -1026 1860 -1021
rect 1865 -1026 1914 -1021
rect 1919 -1026 1966 -1021
rect 871 -1216 1251 -1210
rect 871 -1217 929 -1216
rect 786 -1226 790 -1220
rect 778 -1227 805 -1226
rect 778 -1231 779 -1227
rect 783 -1231 800 -1227
rect 804 -1231 805 -1227
rect 778 -1232 805 -1231
rect 213 -1248 240 -1247
rect 213 -1252 214 -1248
rect 218 -1252 235 -1248
rect 239 -1252 240 -1248
rect 213 -1253 240 -1252
rect 370 -1249 684 -1244
rect 370 -1266 381 -1249
rect 871 -1266 881 -1217
rect 331 -1271 382 -1266
rect 370 -1272 381 -1271
rect 421 -1272 881 -1266
rect 178 -1278 182 -1272
rect -3110 -1288 -3106 -1278
rect 170 -1279 197 -1278
rect 170 -1283 171 -1279
rect 175 -1283 192 -1279
rect 196 -1283 197 -1279
rect 170 -1284 197 -1283
rect 421 -1288 428 -1272
rect -3240 -1293 -3236 -1288
rect -3161 -1292 -3147 -1288
rect -3153 -1293 -3147 -1292
rect -3136 -1293 -3118 -1288
rect -3110 -1293 -3097 -1288
rect -3187 -1304 -3161 -1299
rect -3153 -1307 -3149 -1293
rect -3110 -1296 -3106 -1293
rect -3313 -1347 -3304 -1342
rect -3281 -1343 -3277 -1336
rect -3232 -1343 -3228 -1333
rect -3281 -1348 -3240 -1343
rect -3232 -1348 -3221 -1343
rect 344 -1294 428 -1288
rect 344 -1299 350 -1294
rect 421 -1295 428 -1294
rect 349 -1305 350 -1299
rect 344 -1313 350 -1305
rect 353 -1306 477 -1305
rect 949 -1306 1011 -1305
rect 353 -1310 1012 -1306
rect 353 -1314 358 -1310
rect 452 -1311 1012 -1310
rect 938 -1312 1000 -1311
rect -3118 -1322 -3114 -1316
rect 353 -1322 358 -1319
rect -3126 -1323 -3099 -1322
rect -3126 -1327 -3125 -1323
rect -3121 -1327 -3104 -1323
rect -3100 -1327 -3099 -1323
rect -3126 -1328 -3099 -1327
rect 553 -1345 607 -1342
rect -3281 -1351 -3277 -1348
rect -3232 -1351 -3228 -1348
rect -3296 -1355 -3259 -1351
rect -3296 -1361 -3292 -1355
rect -3263 -1361 -3259 -1355
rect -3161 -1353 -3157 -1347
rect 553 -1349 556 -1345
rect 560 -1349 573 -1345
rect 577 -1349 583 -1345
rect 587 -1349 600 -1345
rect 604 -1349 607 -1345
rect 553 -1351 607 -1349
rect -3169 -1354 -3142 -1353
rect -3169 -1358 -3168 -1354
rect -3164 -1358 -3147 -1354
rect -3143 -1358 -3142 -1354
rect -3169 -1359 -3142 -1358
rect 561 -1356 565 -1351
rect 588 -1356 592 -1351
rect -3240 -1377 -3236 -1371
rect -3248 -1378 -3221 -1377
rect -3304 -1387 -3300 -1381
rect -3271 -1387 -3267 -1381
rect -3248 -1382 -3247 -1378
rect -3243 -1382 -3226 -1378
rect -3222 -1382 -3221 -1378
rect -3248 -1383 -3221 -1382
rect -137 -1380 -73 -1377
rect -137 -1384 -134 -1380
rect -130 -1384 -112 -1380
rect -108 -1384 -102 -1380
rect -98 -1384 -80 -1380
rect -76 -1384 -73 -1380
rect -3312 -1388 -3285 -1387
rect -3312 -1392 -3311 -1388
rect -3307 -1392 -3290 -1388
rect -3286 -1392 -3285 -1388
rect -3312 -1393 -3285 -1392
rect -3279 -1388 -3252 -1387
rect -3279 -1392 -3278 -1388
rect -3274 -1392 -3257 -1388
rect -3253 -1392 -3252 -1388
rect -3279 -1393 -3252 -1392
rect -338 -1388 -150 -1385
rect -137 -1386 -73 -1384
rect -338 -1392 -335 -1388
rect -331 -1392 -313 -1388
rect -309 -1392 -283 -1388
rect -279 -1392 -261 -1388
rect -257 -1392 -231 -1388
rect -227 -1392 -209 -1388
rect -205 -1392 -179 -1388
rect -175 -1392 -157 -1388
rect -153 -1392 -150 -1388
rect -338 -1394 -150 -1392
rect -127 -1392 -123 -1386
rect -95 -1392 -91 -1386
rect -328 -1400 -324 -1394
rect -276 -1400 -272 -1394
rect -224 -1400 -220 -1394
rect -172 -1400 -168 -1394
rect 569 -1416 573 -1396
rect 596 -1416 600 -1396
rect 615 -1415 642 -1412
rect 451 -1420 476 -1419
rect 569 -1420 610 -1416
rect 349 -1421 476 -1420
rect 349 -1425 561 -1421
rect 475 -1426 561 -1425
rect 588 -1430 592 -1420
rect -351 -1449 -328 -1444
rect -351 -1515 -346 -1449
rect -320 -1453 -316 -1440
rect -328 -1457 -316 -1453
rect -298 -1449 -276 -1444
rect -328 -1462 -324 -1457
rect -333 -1511 -328 -1506
rect -320 -1515 -316 -1502
rect -298 -1515 -293 -1449
rect -268 -1453 -264 -1440
rect -216 -1444 -212 -1440
rect -164 -1444 -160 -1440
rect -119 -1444 -115 -1432
rect -87 -1444 -83 -1432
rect -276 -1457 -264 -1453
rect -246 -1449 -224 -1444
rect -216 -1449 -172 -1444
rect -164 -1449 -127 -1444
rect -119 -1449 -95 -1444
rect -87 -1449 -1 -1444
rect -276 -1462 -272 -1457
rect -281 -1511 -276 -1506
rect -268 -1515 -264 -1502
rect -246 -1515 -241 -1449
rect -227 -1472 -224 -1467
rect -216 -1476 -212 -1449
rect -224 -1507 -220 -1496
rect -224 -1511 -212 -1507
rect -351 -1520 -328 -1515
rect -320 -1520 -276 -1515
rect -268 -1520 -224 -1515
rect -320 -1523 -316 -1520
rect -268 -1523 -264 -1520
rect -216 -1523 -212 -1511
rect -194 -1515 -189 -1449
rect -175 -1472 -172 -1467
rect -164 -1476 -160 -1449
rect -119 -1452 -115 -1449
rect -87 -1452 -83 -1449
rect -79 -1450 -1 -1449
rect -127 -1479 -123 -1472
rect -95 -1479 -91 -1472
rect -137 -1481 -73 -1479
rect -137 -1485 -135 -1481
rect -131 -1485 -111 -1481
rect -107 -1485 -103 -1481
rect -99 -1485 -79 -1481
rect -75 -1485 -73 -1481
rect -137 -1487 -73 -1485
rect -172 -1507 -168 -1496
rect -172 -1511 -160 -1507
rect -194 -1520 -172 -1515
rect -164 -1523 -160 -1511
rect -328 -1551 -324 -1543
rect -276 -1551 -272 -1543
rect -224 -1551 -220 -1543
rect -172 -1551 -168 -1543
rect -338 -1552 -150 -1551
rect -338 -1556 -311 -1552
rect -307 -1556 -259 -1552
rect -255 -1556 -207 -1552
rect -203 -1556 -155 -1552
rect -151 -1556 -150 -1552
rect -338 -1557 -150 -1556
rect -345 -1570 -338 -1565
rect -333 -1570 -286 -1565
rect -281 -1570 -232 -1565
rect -227 -1570 -180 -1565
rect -19 -1617 -6 -1450
rect 580 -1476 584 -1470
rect 605 -1476 610 -1420
rect 615 -1419 618 -1415
rect 622 -1419 635 -1415
rect 639 -1419 642 -1415
rect 615 -1421 642 -1419
rect 623 -1426 627 -1421
rect 631 -1476 635 -1466
rect 580 -1480 594 -1476
rect 588 -1481 594 -1480
rect 605 -1481 623 -1476
rect 631 -1477 644 -1476
rect 631 -1481 942 -1477
rect 340 -1487 476 -1486
rect 340 -1491 580 -1487
rect 451 -1492 580 -1491
rect 588 -1495 592 -1481
rect 631 -1484 635 -1481
rect 638 -1482 942 -1481
rect 623 -1510 627 -1504
rect 615 -1511 642 -1510
rect 615 -1515 616 -1511
rect 620 -1515 637 -1511
rect 641 -1515 642 -1511
rect 615 -1516 642 -1515
rect 580 -1541 584 -1535
rect 572 -1542 599 -1541
rect 572 -1546 573 -1542
rect 577 -1546 594 -1542
rect 598 -1546 599 -1542
rect 572 -1547 599 -1546
rect 790 -1575 844 -1572
rect 790 -1579 793 -1575
rect 797 -1579 810 -1575
rect 814 -1579 820 -1575
rect 824 -1579 837 -1575
rect 841 -1579 844 -1575
rect 790 -1581 844 -1579
rect 798 -1586 802 -1581
rect 825 -1586 829 -1581
rect 243 -1598 270 -1595
rect 243 -1602 246 -1598
rect 250 -1602 263 -1598
rect 267 -1602 270 -1598
rect 243 -1604 270 -1602
rect 251 -1609 255 -1604
rect 140 -1617 145 -1615
rect -22 -1622 11 -1617
rect 16 -1622 145 -1617
rect 105 -1626 111 -1625
rect 105 -1630 106 -1626
rect 110 -1630 111 -1626
rect 105 -1633 111 -1630
rect 140 -1633 145 -1622
rect 200 -1628 209 -1625
rect 200 -1632 202 -1628
rect 206 -1632 209 -1628
rect 223 -1632 236 -1629
rect 200 -1633 209 -1632
rect 105 -1637 117 -1633
rect 105 -1647 111 -1637
rect 195 -1637 209 -1633
rect 137 -1645 155 -1641
rect 200 -1645 209 -1637
rect 105 -1651 106 -1647
rect 110 -1651 111 -1647
rect 105 -1652 111 -1651
rect 140 -1655 145 -1645
rect 200 -1649 202 -1645
rect 206 -1649 209 -1645
rect 200 -1652 209 -1649
rect 215 -1655 219 -1652
rect 169 -1659 219 -1655
rect -32 -1664 -16 -1663
rect 169 -1664 173 -1659
rect -32 -1669 173 -1664
rect 223 -1665 227 -1652
rect 230 -1659 236 -1632
rect 554 -1628 608 -1625
rect 935 -1618 942 -1482
rect 1005 -1515 1012 -1311
rect 1072 -1421 1099 -1418
rect 1072 -1425 1075 -1421
rect 1079 -1425 1092 -1421
rect 1096 -1425 1099 -1421
rect 1072 -1427 1099 -1425
rect 1080 -1432 1084 -1427
rect 1005 -1520 1080 -1515
rect 1088 -1524 1092 -1512
rect 1080 -1528 1092 -1524
rect 1080 -1532 1084 -1528
rect 1121 -1558 1148 -1555
rect 1121 -1562 1124 -1558
rect 1128 -1562 1141 -1558
rect 1145 -1562 1148 -1558
rect 1121 -1564 1148 -1562
rect 1129 -1569 1133 -1564
rect 1369 -1574 1396 -1571
rect 1369 -1578 1372 -1574
rect 1376 -1578 1389 -1574
rect 1393 -1578 1396 -1574
rect 1369 -1580 1396 -1578
rect 935 -1623 1065 -1618
rect 1088 -1619 1092 -1612
rect 1137 -1619 1141 -1609
rect 1377 -1585 1381 -1580
rect 935 -1626 942 -1623
rect 1088 -1624 1129 -1619
rect 1137 -1624 1365 -1619
rect 554 -1632 557 -1628
rect 561 -1632 574 -1628
rect 578 -1632 584 -1628
rect 588 -1632 601 -1628
rect 605 -1632 608 -1628
rect 554 -1634 608 -1632
rect 259 -1659 263 -1649
rect 562 -1639 566 -1634
rect 589 -1639 593 -1634
rect 230 -1664 251 -1659
rect 259 -1664 344 -1659
rect 349 -1664 378 -1659
rect -152 -1717 -88 -1714
rect -152 -1721 -149 -1717
rect -145 -1721 -127 -1717
rect -123 -1721 -117 -1717
rect -113 -1721 -95 -1717
rect -91 -1721 -88 -1717
rect -353 -1725 -165 -1722
rect -152 -1723 -88 -1721
rect -353 -1729 -350 -1725
rect -346 -1729 -328 -1725
rect -324 -1729 -298 -1725
rect -294 -1729 -276 -1725
rect -272 -1729 -246 -1725
rect -242 -1729 -224 -1725
rect -220 -1729 -194 -1725
rect -190 -1729 -172 -1725
rect -168 -1729 -165 -1725
rect -353 -1731 -165 -1729
rect -142 -1729 -138 -1723
rect -110 -1729 -106 -1723
rect -343 -1737 -339 -1731
rect -291 -1737 -287 -1731
rect -239 -1737 -235 -1731
rect -187 -1737 -183 -1731
rect -366 -1786 -343 -1781
rect -366 -1852 -361 -1786
rect -335 -1790 -331 -1777
rect -343 -1794 -331 -1790
rect -313 -1786 -291 -1781
rect -343 -1799 -339 -1794
rect -348 -1848 -343 -1843
rect -335 -1852 -331 -1839
rect -313 -1852 -308 -1786
rect -283 -1790 -279 -1777
rect -231 -1781 -227 -1777
rect -179 -1781 -175 -1777
rect -134 -1781 -130 -1769
rect -102 -1781 -98 -1769
rect -32 -1781 -24 -1669
rect -291 -1794 -279 -1790
rect -261 -1786 -239 -1781
rect -231 -1786 -187 -1781
rect -179 -1786 -142 -1781
rect -134 -1786 -110 -1781
rect -102 -1786 -24 -1781
rect -291 -1799 -287 -1794
rect -296 -1848 -291 -1843
rect -283 -1852 -279 -1839
rect -261 -1852 -256 -1786
rect -242 -1809 -239 -1804
rect -231 -1813 -227 -1786
rect -239 -1844 -235 -1833
rect -239 -1848 -227 -1844
rect -366 -1857 -343 -1852
rect -335 -1857 -291 -1852
rect -283 -1857 -239 -1852
rect -335 -1860 -331 -1857
rect -283 -1860 -279 -1857
rect -231 -1860 -227 -1848
rect -209 -1852 -204 -1786
rect -190 -1809 -187 -1804
rect -179 -1813 -175 -1786
rect -134 -1789 -130 -1786
rect -102 -1789 -98 -1786
rect -90 -1788 -24 -1786
rect -32 -1789 -24 -1788
rect -142 -1816 -138 -1809
rect -110 -1816 -106 -1809
rect -152 -1818 -88 -1816
rect -152 -1822 -150 -1818
rect -146 -1822 -126 -1818
rect -122 -1822 -118 -1818
rect -114 -1822 -94 -1818
rect -90 -1822 -88 -1818
rect -152 -1824 -88 -1822
rect -187 -1844 -183 -1833
rect -187 -1848 -175 -1844
rect -209 -1857 -187 -1852
rect -179 -1860 -175 -1848
rect -343 -1888 -339 -1880
rect -291 -1888 -287 -1880
rect -239 -1888 -235 -1880
rect -187 -1888 -183 -1880
rect 66 -1884 71 -1669
rect 105 -1677 111 -1676
rect 105 -1681 106 -1677
rect 110 -1681 111 -1677
rect 105 -1684 111 -1681
rect 140 -1684 145 -1669
rect 200 -1679 209 -1676
rect 200 -1683 202 -1679
rect 206 -1683 209 -1679
rect 200 -1684 209 -1683
rect 105 -1688 117 -1684
rect 105 -1698 111 -1688
rect 195 -1688 209 -1684
rect 137 -1696 155 -1692
rect 200 -1696 209 -1688
rect 105 -1702 106 -1698
rect 110 -1702 111 -1698
rect 105 -1703 111 -1702
rect 140 -1716 145 -1696
rect 200 -1700 202 -1696
rect 206 -1700 209 -1696
rect 200 -1703 209 -1700
rect 259 -1667 263 -1664
rect 215 -1716 219 -1685
rect 806 -1646 810 -1626
rect 833 -1646 837 -1626
rect 1088 -1627 1092 -1624
rect 1137 -1627 1141 -1624
rect 1073 -1631 1110 -1627
rect 1073 -1637 1077 -1631
rect 1106 -1637 1110 -1631
rect 852 -1645 879 -1642
rect 806 -1650 847 -1646
rect 791 -1652 798 -1651
rect 251 -1693 255 -1687
rect 243 -1694 270 -1693
rect 243 -1698 244 -1694
rect 248 -1698 265 -1694
rect 269 -1698 270 -1694
rect 243 -1699 270 -1698
rect 570 -1699 574 -1679
rect 597 -1699 601 -1679
rect 730 -1656 798 -1652
rect 730 -1657 796 -1656
rect 616 -1698 643 -1695
rect 570 -1703 611 -1699
rect 349 -1704 478 -1703
rect 349 -1708 562 -1704
rect 453 -1709 562 -1708
rect 589 -1713 593 -1703
rect 140 -1719 219 -1716
rect 160 -1742 214 -1739
rect 160 -1746 163 -1742
rect 167 -1746 180 -1742
rect 184 -1746 190 -1742
rect 194 -1746 207 -1742
rect 211 -1746 214 -1742
rect 160 -1748 214 -1746
rect 168 -1753 172 -1748
rect 195 -1753 199 -1748
rect 581 -1759 585 -1753
rect 606 -1759 611 -1703
rect 616 -1702 619 -1698
rect 623 -1702 636 -1698
rect 640 -1702 643 -1698
rect 616 -1704 643 -1702
rect 624 -1709 628 -1704
rect 632 -1759 636 -1749
rect 730 -1759 735 -1657
rect 825 -1660 829 -1650
rect 817 -1706 821 -1700
rect 842 -1706 847 -1650
rect 852 -1649 855 -1645
rect 859 -1649 872 -1645
rect 876 -1649 879 -1645
rect 852 -1651 879 -1649
rect 860 -1656 864 -1651
rect 1129 -1653 1133 -1647
rect 1121 -1654 1148 -1653
rect 1065 -1663 1069 -1657
rect 1098 -1663 1102 -1657
rect 1121 -1658 1122 -1654
rect 1126 -1658 1143 -1654
rect 1147 -1658 1148 -1654
rect 1121 -1659 1148 -1658
rect 1057 -1664 1084 -1663
rect 1057 -1668 1058 -1664
rect 1062 -1668 1079 -1664
rect 1083 -1668 1084 -1664
rect 1057 -1669 1084 -1668
rect 1090 -1664 1117 -1663
rect 1090 -1668 1091 -1664
rect 1095 -1668 1112 -1664
rect 1116 -1668 1117 -1664
rect 1090 -1669 1117 -1668
rect 1360 -1668 1365 -1624
rect 2198 -1586 2262 -1583
rect 2198 -1590 2201 -1586
rect 2205 -1590 2223 -1586
rect 2227 -1590 2233 -1586
rect 2237 -1590 2255 -1586
rect 2259 -1590 2262 -1586
rect 1997 -1594 2185 -1591
rect 2198 -1592 2262 -1590
rect 1997 -1598 2000 -1594
rect 2004 -1598 2022 -1594
rect 2026 -1598 2052 -1594
rect 2056 -1598 2074 -1594
rect 2078 -1598 2104 -1594
rect 2108 -1598 2126 -1594
rect 2130 -1598 2156 -1594
rect 2160 -1598 2178 -1594
rect 2182 -1598 2185 -1594
rect 1997 -1600 2185 -1598
rect 2208 -1598 2212 -1592
rect 2240 -1598 2244 -1592
rect 2007 -1606 2011 -1600
rect 2059 -1606 2063 -1600
rect 2111 -1606 2115 -1600
rect 2163 -1606 2167 -1600
rect 1787 -1639 1814 -1636
rect 1787 -1643 1790 -1639
rect 1794 -1643 1807 -1639
rect 1811 -1643 1814 -1639
rect 1787 -1645 1814 -1643
rect 1795 -1650 1799 -1645
rect 1559 -1656 1654 -1655
rect 1360 -1673 1377 -1668
rect 1385 -1677 1389 -1665
rect 868 -1706 872 -1696
rect 1377 -1681 1389 -1677
rect 1448 -1658 1654 -1656
rect 1684 -1658 1689 -1656
rect 1448 -1660 1689 -1658
rect 1377 -1685 1381 -1681
rect 817 -1710 831 -1706
rect 825 -1711 831 -1710
rect 842 -1711 860 -1706
rect 868 -1707 881 -1706
rect 868 -1711 1017 -1707
rect 581 -1763 595 -1759
rect 589 -1764 595 -1763
rect 606 -1764 624 -1759
rect 632 -1764 735 -1759
rect 751 -1722 817 -1717
rect 331 -1770 455 -1769
rect 331 -1774 581 -1770
rect 453 -1775 581 -1774
rect 453 -1776 478 -1775
rect 589 -1778 593 -1764
rect 632 -1767 636 -1764
rect 176 -1813 180 -1793
rect 203 -1813 207 -1793
rect 222 -1812 249 -1809
rect 176 -1817 217 -1813
rect 104 -1823 168 -1818
rect 195 -1827 199 -1817
rect 187 -1873 191 -1867
rect 212 -1873 217 -1817
rect 222 -1816 225 -1812
rect 229 -1816 242 -1812
rect 246 -1816 249 -1812
rect 222 -1818 249 -1816
rect 624 -1793 628 -1787
rect 616 -1794 643 -1793
rect 616 -1798 617 -1794
rect 621 -1798 638 -1794
rect 642 -1798 643 -1794
rect 616 -1799 643 -1798
rect 230 -1823 234 -1818
rect 581 -1824 585 -1818
rect 573 -1825 600 -1824
rect 573 -1829 574 -1825
rect 578 -1829 595 -1825
rect 599 -1829 600 -1825
rect 573 -1830 600 -1829
rect 453 -1840 478 -1838
rect 322 -1841 478 -1840
rect 751 -1841 756 -1722
rect 825 -1725 829 -1711
rect 868 -1714 872 -1711
rect 875 -1712 1017 -1711
rect 860 -1740 864 -1734
rect 852 -1741 879 -1740
rect 852 -1745 853 -1741
rect 857 -1745 874 -1741
rect 878 -1745 879 -1741
rect 852 -1746 879 -1745
rect 817 -1771 821 -1765
rect 809 -1772 836 -1771
rect 809 -1776 810 -1772
rect 814 -1776 831 -1772
rect 835 -1776 836 -1772
rect 809 -1777 836 -1776
rect 799 -1786 853 -1783
rect 799 -1790 802 -1786
rect 806 -1790 819 -1786
rect 823 -1790 829 -1786
rect 833 -1790 846 -1786
rect 850 -1790 853 -1786
rect 799 -1792 853 -1790
rect 807 -1797 811 -1792
rect 834 -1797 838 -1792
rect 1008 -1815 1017 -1712
rect 1083 -1721 1110 -1718
rect 1083 -1725 1086 -1721
rect 1090 -1725 1103 -1721
rect 1107 -1725 1110 -1721
rect 1083 -1727 1110 -1725
rect 1091 -1732 1095 -1727
rect 1418 -1711 1445 -1708
rect 1418 -1715 1421 -1711
rect 1425 -1715 1438 -1711
rect 1442 -1715 1445 -1711
rect 1418 -1717 1445 -1715
rect 1426 -1722 1430 -1717
rect 1008 -1820 1091 -1815
rect 1099 -1824 1103 -1812
rect 322 -1845 756 -1841
rect 475 -1846 756 -1845
rect 815 -1857 819 -1837
rect 842 -1857 846 -1837
rect 1091 -1828 1103 -1824
rect 1334 -1776 1362 -1771
rect 1385 -1772 1389 -1765
rect 1434 -1772 1438 -1762
rect 1448 -1772 1452 -1660
rect 1649 -1663 1689 -1660
rect 1649 -1667 1655 -1666
rect 1649 -1671 1650 -1667
rect 1654 -1671 1655 -1667
rect 1649 -1674 1655 -1671
rect 1684 -1674 1689 -1663
rect 1744 -1669 1753 -1666
rect 1744 -1673 1746 -1669
rect 1750 -1673 1753 -1669
rect 1767 -1673 1780 -1670
rect 1744 -1674 1753 -1673
rect 1649 -1678 1661 -1674
rect 1649 -1688 1655 -1678
rect 1739 -1678 1753 -1674
rect 1681 -1686 1699 -1682
rect 1744 -1686 1753 -1678
rect 1649 -1692 1650 -1688
rect 1654 -1692 1655 -1688
rect 1649 -1693 1655 -1692
rect 1684 -1696 1689 -1686
rect 1744 -1690 1746 -1686
rect 1750 -1690 1753 -1686
rect 1744 -1693 1753 -1690
rect 1759 -1696 1763 -1693
rect 1713 -1700 1763 -1696
rect 1713 -1705 1717 -1700
rect 1091 -1832 1095 -1828
rect 861 -1856 888 -1853
rect 815 -1861 856 -1857
rect 800 -1863 807 -1862
rect 238 -1873 242 -1863
rect 736 -1867 807 -1863
rect 736 -1868 803 -1867
rect 187 -1877 201 -1873
rect 195 -1878 201 -1877
rect 212 -1878 230 -1873
rect 238 -1878 353 -1873
rect 358 -1878 391 -1873
rect -353 -1889 -165 -1888
rect 66 -1889 187 -1884
rect -353 -1893 -326 -1889
rect -322 -1893 -274 -1889
rect -270 -1893 -222 -1889
rect -218 -1893 -170 -1889
rect -166 -1893 -165 -1889
rect 195 -1892 199 -1878
rect 238 -1881 242 -1878
rect -353 -1894 -165 -1893
rect -360 -1907 -353 -1902
rect -348 -1907 -301 -1902
rect -296 -1907 -247 -1902
rect -242 -1907 -195 -1902
rect 550 -1899 604 -1896
rect 230 -1907 234 -1901
rect 550 -1903 553 -1899
rect 557 -1903 570 -1899
rect 574 -1903 580 -1899
rect 584 -1903 597 -1899
rect 601 -1903 604 -1899
rect 550 -1905 604 -1903
rect 222 -1908 249 -1907
rect 222 -1912 223 -1908
rect 227 -1912 244 -1908
rect 248 -1912 249 -1908
rect 222 -1913 249 -1912
rect 558 -1910 562 -1905
rect 585 -1910 589 -1905
rect 187 -1938 191 -1932
rect 179 -1939 206 -1938
rect 179 -1943 180 -1939
rect 184 -1943 201 -1939
rect 205 -1943 206 -1939
rect 179 -1944 206 -1943
rect 566 -1970 570 -1950
rect 593 -1970 597 -1950
rect 612 -1969 639 -1966
rect 566 -1974 607 -1970
rect 304 -1975 478 -1974
rect 304 -1979 558 -1975
rect 453 -1980 558 -1979
rect 585 -1984 589 -1974
rect 577 -2030 581 -2024
rect 602 -2030 607 -1974
rect 612 -1973 615 -1969
rect 619 -1973 632 -1969
rect 636 -1973 639 -1969
rect 612 -1975 639 -1973
rect 620 -1980 624 -1975
rect 628 -2030 632 -2020
rect 736 -2030 741 -1868
rect 834 -1871 838 -1861
rect 826 -1917 830 -1911
rect 851 -1917 856 -1861
rect 861 -1860 864 -1856
rect 868 -1860 881 -1856
rect 885 -1860 888 -1856
rect 861 -1862 888 -1860
rect 869 -1867 873 -1862
rect 877 -1917 881 -1907
rect 1132 -1858 1159 -1855
rect 1132 -1862 1135 -1858
rect 1139 -1862 1152 -1858
rect 1156 -1862 1159 -1858
rect 1132 -1864 1159 -1862
rect 1140 -1869 1144 -1864
rect 826 -1921 840 -1917
rect 834 -1922 840 -1921
rect 851 -1922 869 -1917
rect 877 -1918 1014 -1917
rect 877 -1922 1076 -1918
rect 800 -1929 826 -1928
rect 577 -2034 591 -2030
rect 585 -2035 591 -2034
rect 602 -2035 620 -2030
rect 628 -2035 741 -2030
rect 775 -1933 826 -1929
rect 775 -1934 816 -1933
rect 307 -2045 308 -2040
rect 313 -2041 455 -2040
rect 313 -2045 577 -2041
rect 452 -2046 577 -2045
rect 452 -2047 477 -2046
rect 585 -2049 589 -2035
rect 628 -2038 632 -2035
rect 620 -2064 624 -2058
rect 612 -2065 639 -2064
rect 612 -2069 613 -2065
rect 617 -2069 634 -2065
rect 638 -2069 639 -2065
rect 612 -2070 639 -2069
rect 775 -2073 780 -1934
rect 834 -1936 838 -1922
rect 877 -1925 881 -1922
rect 907 -1923 1076 -1922
rect 1099 -1919 1103 -1912
rect 1148 -1919 1152 -1909
rect 1334 -1919 1339 -1776
rect 1385 -1777 1426 -1772
rect 1434 -1777 1452 -1772
rect 1385 -1780 1389 -1777
rect 1434 -1780 1438 -1777
rect 1448 -1779 1452 -1777
rect 1563 -1710 1717 -1705
rect 1767 -1706 1771 -1693
rect 1774 -1700 1780 -1673
rect 1803 -1700 1807 -1690
rect 1984 -1655 2007 -1650
rect 1984 -1700 1989 -1655
rect 2015 -1659 2019 -1646
rect 1774 -1705 1795 -1700
rect 1803 -1705 1989 -1700
rect 1370 -1784 1407 -1780
rect 1370 -1790 1374 -1784
rect 1403 -1790 1407 -1784
rect 1426 -1806 1430 -1800
rect 1418 -1807 1445 -1806
rect 1362 -1816 1366 -1810
rect 1395 -1816 1399 -1810
rect 1418 -1811 1419 -1807
rect 1423 -1811 1440 -1807
rect 1444 -1811 1445 -1807
rect 1418 -1812 1445 -1811
rect 1354 -1817 1381 -1816
rect 1354 -1821 1355 -1817
rect 1359 -1821 1376 -1817
rect 1380 -1821 1381 -1817
rect 1354 -1822 1381 -1821
rect 1387 -1817 1414 -1816
rect 1387 -1821 1388 -1817
rect 1392 -1821 1409 -1817
rect 1413 -1821 1414 -1817
rect 1387 -1822 1414 -1821
rect 1099 -1924 1140 -1919
rect 1148 -1924 1339 -1919
rect 1375 -1860 1380 -1858
rect 1563 -1860 1568 -1710
rect 1649 -1718 1655 -1717
rect 1649 -1722 1650 -1718
rect 1654 -1722 1655 -1718
rect 1649 -1725 1655 -1722
rect 1684 -1725 1689 -1710
rect 1744 -1720 1753 -1717
rect 1744 -1724 1746 -1720
rect 1750 -1724 1753 -1720
rect 1744 -1725 1753 -1724
rect 1649 -1729 1661 -1725
rect 1649 -1739 1655 -1729
rect 1739 -1729 1753 -1725
rect 1681 -1737 1699 -1733
rect 1744 -1737 1753 -1729
rect 1649 -1743 1650 -1739
rect 1654 -1743 1655 -1739
rect 1649 -1744 1655 -1743
rect 1684 -1757 1689 -1737
rect 1744 -1741 1746 -1737
rect 1750 -1741 1753 -1737
rect 1744 -1744 1753 -1741
rect 1803 -1708 1807 -1705
rect 1812 -1708 1989 -1705
rect 2007 -1663 2019 -1659
rect 2037 -1655 2059 -1650
rect 2007 -1668 2011 -1663
rect 1759 -1757 1763 -1726
rect 1984 -1721 1989 -1708
rect 2002 -1717 2007 -1712
rect 2015 -1721 2019 -1708
rect 2037 -1721 2042 -1655
rect 2067 -1659 2071 -1646
rect 2119 -1650 2123 -1646
rect 2171 -1650 2175 -1646
rect 2216 -1650 2220 -1638
rect 2248 -1650 2252 -1638
rect 2059 -1663 2071 -1659
rect 2089 -1655 2111 -1650
rect 2119 -1655 2163 -1650
rect 2171 -1655 2208 -1650
rect 2216 -1655 2240 -1650
rect 2248 -1655 2262 -1650
rect 2059 -1668 2063 -1663
rect 2054 -1717 2059 -1712
rect 2067 -1721 2071 -1708
rect 2089 -1721 2094 -1655
rect 2108 -1678 2111 -1673
rect 2119 -1682 2123 -1655
rect 2111 -1713 2115 -1702
rect 2111 -1717 2123 -1713
rect 1984 -1726 2007 -1721
rect 2015 -1726 2059 -1721
rect 2067 -1726 2111 -1721
rect 1795 -1734 1799 -1728
rect 2015 -1729 2019 -1726
rect 2067 -1729 2071 -1726
rect 2119 -1729 2123 -1717
rect 2141 -1721 2146 -1655
rect 2160 -1678 2163 -1673
rect 2171 -1682 2175 -1655
rect 2216 -1658 2220 -1655
rect 2248 -1658 2252 -1655
rect 2208 -1685 2212 -1678
rect 2240 -1685 2244 -1678
rect 2198 -1687 2262 -1685
rect 2198 -1691 2200 -1687
rect 2204 -1691 2224 -1687
rect 2228 -1691 2232 -1687
rect 2236 -1691 2256 -1687
rect 2260 -1691 2262 -1687
rect 2198 -1693 2262 -1691
rect 2163 -1713 2167 -1702
rect 2163 -1717 2175 -1713
rect 2141 -1726 2163 -1721
rect 2171 -1729 2175 -1717
rect 1787 -1735 1814 -1734
rect 1787 -1739 1788 -1735
rect 1792 -1739 1809 -1735
rect 1813 -1739 1814 -1735
rect 1787 -1740 1814 -1739
rect 2007 -1757 2011 -1749
rect 2059 -1757 2063 -1749
rect 2111 -1757 2115 -1749
rect 2163 -1757 2167 -1749
rect 1684 -1760 1763 -1757
rect 1997 -1758 2185 -1757
rect 1997 -1762 2024 -1758
rect 2028 -1762 2076 -1758
rect 2080 -1762 2128 -1758
rect 2132 -1762 2180 -1758
rect 2184 -1762 2185 -1758
rect 1997 -1763 2185 -1762
rect 1990 -1776 1997 -1771
rect 2002 -1776 2049 -1771
rect 2054 -1776 2103 -1771
rect 2108 -1776 2155 -1771
rect 1375 -1868 1568 -1860
rect 1099 -1927 1103 -1924
rect 1148 -1927 1152 -1924
rect 1084 -1931 1121 -1927
rect 1084 -1937 1088 -1931
rect 1117 -1937 1121 -1931
rect 869 -1951 873 -1945
rect 861 -1952 888 -1951
rect 861 -1956 862 -1952
rect 866 -1956 883 -1952
rect 887 -1956 888 -1952
rect 861 -1957 888 -1956
rect 1140 -1953 1144 -1947
rect 1132 -1954 1159 -1953
rect 1076 -1963 1080 -1957
rect 1109 -1963 1113 -1957
rect 1132 -1958 1133 -1954
rect 1137 -1958 1154 -1954
rect 1158 -1958 1159 -1954
rect 1132 -1959 1159 -1958
rect 1068 -1964 1095 -1963
rect 1068 -1968 1069 -1964
rect 1073 -1968 1090 -1964
rect 1094 -1968 1095 -1964
rect 1068 -1969 1095 -1968
rect 1101 -1964 1128 -1963
rect 1101 -1968 1102 -1964
rect 1106 -1968 1123 -1964
rect 1127 -1968 1128 -1964
rect 1101 -1969 1128 -1968
rect 826 -1982 830 -1976
rect 818 -1983 845 -1982
rect 818 -1987 819 -1983
rect 823 -1987 840 -1983
rect 844 -1987 845 -1983
rect 818 -1988 845 -1987
rect 1375 -2048 1380 -1868
rect 1563 -1870 1568 -1868
rect 690 -2082 780 -2073
rect 1010 -2053 1381 -2048
rect 690 -2088 703 -2082
rect 577 -2095 581 -2089
rect 569 -2096 596 -2095
rect 569 -2100 570 -2096
rect 574 -2100 591 -2096
rect 595 -2100 596 -2096
rect 569 -2101 596 -2100
rect 538 -2148 592 -2145
rect 538 -2152 541 -2148
rect 545 -2152 558 -2148
rect 562 -2152 568 -2148
rect 572 -2152 585 -2148
rect 589 -2152 592 -2148
rect 538 -2154 592 -2152
rect 546 -2159 550 -2154
rect 573 -2159 577 -2154
rect 554 -2219 558 -2199
rect 581 -2219 585 -2199
rect 600 -2218 627 -2215
rect 554 -2223 595 -2219
rect 343 -2228 344 -2223
rect 349 -2224 476 -2223
rect 349 -2228 546 -2224
rect 451 -2229 546 -2228
rect 573 -2233 577 -2223
rect 565 -2279 569 -2273
rect 590 -2279 595 -2223
rect 600 -2222 603 -2218
rect 607 -2222 620 -2218
rect 624 -2222 627 -2218
rect 600 -2224 627 -2222
rect 608 -2229 612 -2224
rect 616 -2279 620 -2269
rect 690 -2279 702 -2088
rect 1010 -2099 1017 -2053
rect 803 -2104 1018 -2099
rect 565 -2283 579 -2279
rect 573 -2284 579 -2283
rect 590 -2284 608 -2279
rect 616 -2284 703 -2279
rect 331 -2290 455 -2289
rect 331 -2294 565 -2290
rect 453 -2295 565 -2294
rect 453 -2296 478 -2295
rect 573 -2298 577 -2284
rect 616 -2287 620 -2284
rect 690 -2287 702 -2284
rect -152 -2324 -88 -2321
rect -152 -2328 -149 -2324
rect -145 -2328 -127 -2324
rect -123 -2328 -117 -2324
rect -113 -2328 -95 -2324
rect -91 -2328 -88 -2324
rect -353 -2332 -165 -2329
rect -152 -2330 -88 -2328
rect -353 -2336 -350 -2332
rect -346 -2336 -328 -2332
rect -324 -2336 -298 -2332
rect -294 -2336 -276 -2332
rect -272 -2336 -246 -2332
rect -242 -2336 -224 -2332
rect -220 -2336 -194 -2332
rect -190 -2336 -172 -2332
rect -168 -2336 -165 -2332
rect -353 -2338 -165 -2336
rect -142 -2336 -138 -2330
rect -110 -2336 -106 -2330
rect -343 -2344 -339 -2338
rect -291 -2344 -287 -2338
rect -239 -2344 -235 -2338
rect -187 -2344 -183 -2338
rect 608 -2313 612 -2307
rect 600 -2314 627 -2313
rect 600 -2318 601 -2314
rect 605 -2318 622 -2314
rect 626 -2318 627 -2314
rect 600 -2319 627 -2318
rect 565 -2344 569 -2338
rect 557 -2345 584 -2344
rect 557 -2349 558 -2345
rect 562 -2349 579 -2345
rect 583 -2349 584 -2345
rect 557 -2350 584 -2349
rect -366 -2393 -343 -2388
rect -366 -2459 -361 -2393
rect -335 -2397 -331 -2384
rect -343 -2401 -331 -2397
rect -313 -2393 -291 -2388
rect -343 -2406 -339 -2401
rect -348 -2455 -343 -2450
rect -335 -2459 -331 -2446
rect -313 -2459 -308 -2393
rect -283 -2397 -279 -2384
rect -231 -2388 -227 -2384
rect -179 -2388 -175 -2384
rect -134 -2388 -130 -2376
rect -102 -2388 -98 -2376
rect 360 -2383 362 -2378
rect 367 -2379 478 -2378
rect 803 -2379 808 -2104
rect 911 -2105 1018 -2104
rect 367 -2383 808 -2379
rect 453 -2384 808 -2383
rect -93 -2388 -19 -2387
rect -291 -2401 -279 -2397
rect -261 -2393 -239 -2388
rect -231 -2393 -187 -2388
rect -179 -2393 -142 -2388
rect -134 -2393 -110 -2388
rect -102 -2393 -19 -2388
rect -291 -2406 -287 -2401
rect -296 -2455 -291 -2450
rect -283 -2459 -279 -2446
rect -261 -2459 -256 -2393
rect -242 -2416 -239 -2411
rect -231 -2420 -227 -2393
rect -239 -2451 -235 -2440
rect -239 -2455 -227 -2451
rect -366 -2464 -343 -2459
rect -335 -2464 -291 -2459
rect -283 -2464 -239 -2459
rect -335 -2467 -331 -2464
rect -283 -2467 -279 -2464
rect -231 -2467 -227 -2455
rect -209 -2459 -204 -2393
rect -190 -2416 -187 -2411
rect -179 -2420 -175 -2393
rect -134 -2396 -130 -2393
rect -102 -2396 -98 -2393
rect -142 -2423 -138 -2416
rect -110 -2423 -106 -2416
rect -152 -2425 -88 -2423
rect -152 -2429 -150 -2425
rect -146 -2429 -126 -2425
rect -122 -2429 -118 -2425
rect -114 -2429 -94 -2425
rect -90 -2429 -88 -2425
rect -152 -2431 -88 -2429
rect -187 -2451 -183 -2440
rect -187 -2455 -175 -2451
rect -209 -2464 -187 -2459
rect -179 -2467 -175 -2455
rect -343 -2495 -339 -2487
rect -291 -2495 -287 -2487
rect -239 -2495 -235 -2487
rect -187 -2495 -183 -2487
rect -29 -2492 -19 -2393
rect 568 -2455 1248 -2454
rect 523 -2459 1248 -2455
rect 523 -2460 571 -2459
rect 240 -2473 267 -2470
rect 240 -2477 243 -2473
rect 247 -2477 260 -2473
rect 264 -2477 267 -2473
rect 240 -2479 267 -2477
rect 248 -2484 252 -2479
rect 137 -2492 142 -2490
rect -353 -2496 -165 -2495
rect -353 -2500 -326 -2496
rect -322 -2500 -274 -2496
rect -270 -2500 -222 -2496
rect -218 -2500 -170 -2496
rect -166 -2500 -165 -2496
rect -29 -2497 8 -2492
rect 13 -2497 142 -2492
rect -29 -2498 -19 -2497
rect -353 -2501 -165 -2500
rect 102 -2501 108 -2500
rect 102 -2505 103 -2501
rect 107 -2505 108 -2501
rect 102 -2508 108 -2505
rect 137 -2508 142 -2497
rect 197 -2503 206 -2500
rect 197 -2507 199 -2503
rect 203 -2507 206 -2503
rect 220 -2507 233 -2504
rect 197 -2508 206 -2507
rect -360 -2514 -353 -2509
rect -348 -2514 -301 -2509
rect -296 -2514 -247 -2509
rect -242 -2514 -195 -2509
rect 102 -2512 114 -2508
rect 102 -2522 108 -2512
rect 192 -2512 206 -2508
rect 134 -2520 152 -2516
rect 197 -2520 206 -2512
rect 102 -2526 103 -2522
rect 107 -2526 108 -2522
rect 102 -2527 108 -2526
rect 137 -2530 142 -2520
rect 197 -2524 199 -2520
rect 203 -2524 206 -2520
rect 197 -2527 206 -2524
rect 212 -2530 216 -2527
rect 166 -2534 216 -2530
rect 166 -2539 170 -2534
rect -26 -2544 170 -2539
rect 220 -2540 224 -2527
rect 227 -2534 233 -2507
rect 256 -2534 260 -2524
rect 227 -2539 248 -2534
rect 256 -2539 362 -2534
rect 367 -2539 387 -2534
rect -152 -2594 -88 -2591
rect -152 -2598 -149 -2594
rect -145 -2598 -127 -2594
rect -123 -2598 -117 -2594
rect -113 -2598 -95 -2594
rect -91 -2598 -88 -2594
rect -353 -2602 -165 -2599
rect -152 -2600 -88 -2598
rect -353 -2606 -350 -2602
rect -346 -2606 -328 -2602
rect -324 -2606 -298 -2602
rect -294 -2606 -276 -2602
rect -272 -2606 -246 -2602
rect -242 -2606 -224 -2602
rect -220 -2606 -194 -2602
rect -190 -2606 -172 -2602
rect -168 -2606 -165 -2602
rect -353 -2608 -165 -2606
rect -142 -2606 -138 -2600
rect -110 -2606 -106 -2600
rect -343 -2614 -339 -2608
rect -291 -2614 -287 -2608
rect -239 -2614 -235 -2608
rect -187 -2614 -183 -2608
rect -366 -2663 -343 -2658
rect -366 -2729 -361 -2663
rect -335 -2667 -331 -2654
rect -343 -2671 -331 -2667
rect -313 -2663 -291 -2658
rect -343 -2676 -339 -2671
rect -348 -2725 -343 -2720
rect -335 -2729 -331 -2716
rect -313 -2729 -308 -2663
rect -283 -2667 -279 -2654
rect -231 -2658 -227 -2654
rect -179 -2658 -175 -2654
rect -134 -2658 -130 -2646
rect -102 -2658 -98 -2646
rect -26 -2658 -20 -2544
rect -291 -2671 -279 -2667
rect -261 -2663 -239 -2658
rect -231 -2663 -187 -2658
rect -179 -2663 -142 -2658
rect -134 -2663 -110 -2658
rect -102 -2663 -20 -2658
rect -291 -2676 -287 -2671
rect -296 -2725 -291 -2720
rect -283 -2729 -279 -2716
rect -261 -2729 -256 -2663
rect -242 -2686 -239 -2681
rect -231 -2690 -227 -2663
rect -239 -2721 -235 -2710
rect -239 -2725 -227 -2721
rect -366 -2734 -343 -2729
rect -335 -2734 -291 -2729
rect -283 -2734 -239 -2729
rect -335 -2737 -331 -2734
rect -283 -2737 -279 -2734
rect -231 -2737 -227 -2725
rect -209 -2729 -204 -2663
rect -190 -2686 -187 -2681
rect -179 -2690 -175 -2663
rect -134 -2666 -130 -2663
rect -102 -2666 -98 -2663
rect -142 -2693 -138 -2686
rect -110 -2693 -106 -2686
rect -152 -2695 -88 -2693
rect -152 -2699 -150 -2695
rect -146 -2699 -126 -2695
rect -122 -2699 -118 -2695
rect -114 -2699 -94 -2695
rect -90 -2699 -88 -2695
rect -152 -2701 -88 -2699
rect -187 -2721 -183 -2710
rect -187 -2725 -175 -2721
rect -209 -2734 -187 -2729
rect -179 -2737 -175 -2725
rect -343 -2765 -339 -2757
rect -291 -2765 -287 -2757
rect -239 -2765 -235 -2757
rect -187 -2765 -183 -2757
rect 63 -2759 68 -2544
rect 102 -2552 108 -2551
rect 102 -2556 103 -2552
rect 107 -2556 108 -2552
rect 102 -2559 108 -2556
rect 137 -2559 142 -2544
rect 197 -2554 206 -2551
rect 197 -2558 199 -2554
rect 203 -2558 206 -2554
rect 197 -2559 206 -2558
rect 102 -2563 114 -2559
rect 102 -2573 108 -2563
rect 192 -2563 206 -2559
rect 134 -2571 152 -2567
rect 197 -2571 206 -2563
rect 102 -2577 103 -2573
rect 107 -2577 108 -2573
rect 102 -2578 108 -2577
rect 137 -2591 142 -2571
rect 197 -2575 199 -2571
rect 203 -2575 206 -2571
rect 197 -2578 206 -2575
rect 256 -2542 260 -2539
rect 212 -2591 216 -2560
rect 248 -2568 252 -2562
rect 240 -2569 267 -2568
rect 240 -2573 241 -2569
rect 245 -2573 262 -2569
rect 266 -2573 267 -2569
rect 240 -2574 267 -2573
rect 137 -2594 216 -2591
rect 157 -2617 211 -2614
rect 157 -2621 160 -2617
rect 164 -2621 177 -2617
rect 181 -2621 187 -2617
rect 191 -2621 204 -2617
rect 208 -2621 211 -2617
rect 157 -2623 211 -2621
rect 165 -2628 169 -2623
rect 192 -2628 196 -2623
rect 173 -2688 177 -2668
rect 200 -2688 204 -2668
rect 219 -2687 246 -2684
rect 173 -2692 214 -2688
rect 101 -2698 165 -2693
rect 192 -2702 196 -2692
rect 184 -2748 188 -2742
rect 209 -2748 214 -2692
rect 219 -2691 222 -2687
rect 226 -2691 239 -2687
rect 243 -2691 246 -2687
rect 219 -2693 246 -2691
rect 227 -2698 231 -2693
rect 235 -2748 239 -2738
rect 523 -2748 528 -2460
rect 850 -2490 1218 -2485
rect 631 -2495 685 -2492
rect 631 -2499 634 -2495
rect 638 -2499 651 -2495
rect 655 -2499 661 -2495
rect 665 -2499 678 -2495
rect 682 -2499 685 -2495
rect 631 -2501 685 -2499
rect 639 -2506 643 -2501
rect 666 -2506 670 -2501
rect 647 -2566 651 -2546
rect 674 -2566 678 -2546
rect 693 -2565 720 -2562
rect 647 -2570 688 -2566
rect 568 -2572 639 -2571
rect 184 -2752 198 -2748
rect 192 -2753 198 -2752
rect 209 -2753 227 -2748
rect 235 -2753 528 -2748
rect 537 -2576 639 -2572
rect 537 -2577 571 -2576
rect 63 -2764 184 -2759
rect -353 -2766 -165 -2765
rect -353 -2770 -326 -2766
rect -322 -2770 -274 -2766
rect -270 -2770 -222 -2766
rect -218 -2770 -170 -2766
rect -166 -2770 -165 -2766
rect 192 -2767 196 -2753
rect 235 -2756 239 -2753
rect -353 -2771 -165 -2770
rect -360 -2784 -353 -2779
rect -348 -2784 -301 -2779
rect -296 -2784 -247 -2779
rect -242 -2784 -195 -2779
rect 537 -2765 542 -2577
rect 666 -2580 670 -2570
rect 658 -2626 662 -2620
rect 683 -2626 688 -2570
rect 693 -2569 696 -2565
rect 700 -2569 713 -2565
rect 717 -2569 720 -2565
rect 693 -2571 720 -2569
rect 701 -2576 705 -2571
rect 709 -2626 713 -2616
rect 850 -2626 855 -2490
rect 966 -2547 1020 -2544
rect 966 -2551 969 -2547
rect 973 -2551 986 -2547
rect 990 -2551 996 -2547
rect 1000 -2551 1013 -2547
rect 1017 -2551 1020 -2547
rect 966 -2553 1020 -2551
rect 974 -2558 978 -2553
rect 1001 -2558 1005 -2553
rect 982 -2618 986 -2598
rect 1009 -2618 1013 -2598
rect 1028 -2617 1055 -2614
rect 982 -2622 1023 -2618
rect 658 -2630 672 -2626
rect 666 -2631 672 -2630
rect 683 -2631 701 -2626
rect 709 -2631 855 -2626
rect 963 -2628 974 -2623
rect 568 -2638 658 -2637
rect 352 -2770 353 -2765
rect 358 -2770 542 -2765
rect 550 -2642 658 -2638
rect 550 -2643 571 -2642
rect 550 -2774 555 -2643
rect 666 -2645 670 -2631
rect 709 -2634 713 -2631
rect 963 -2641 971 -2628
rect 1001 -2632 1005 -2622
rect 902 -2643 971 -2641
rect 855 -2648 971 -2643
rect 701 -2660 705 -2654
rect 693 -2661 720 -2660
rect 693 -2665 694 -2661
rect 698 -2665 715 -2661
rect 719 -2665 720 -2661
rect 693 -2666 720 -2665
rect 658 -2691 662 -2685
rect 650 -2692 677 -2691
rect 650 -2696 651 -2692
rect 655 -2696 672 -2692
rect 676 -2696 677 -2692
rect 650 -2697 677 -2696
rect 227 -2782 231 -2776
rect 367 -2779 555 -2774
rect 632 -2778 686 -2775
rect 632 -2782 635 -2778
rect 639 -2782 652 -2778
rect 656 -2782 662 -2778
rect 666 -2782 679 -2778
rect 683 -2782 686 -2778
rect 219 -2783 246 -2782
rect 219 -2787 220 -2783
rect 224 -2787 241 -2783
rect 245 -2787 246 -2783
rect 632 -2784 686 -2782
rect 219 -2788 246 -2787
rect 640 -2789 644 -2784
rect 667 -2789 671 -2784
rect 184 -2813 188 -2807
rect 176 -2814 203 -2813
rect 176 -2818 177 -2814
rect 181 -2818 198 -2814
rect 202 -2818 203 -2814
rect 176 -2819 203 -2818
rect 648 -2849 652 -2829
rect 675 -2849 679 -2829
rect 694 -2848 721 -2845
rect 648 -2853 689 -2849
rect 568 -2855 640 -2854
rect 361 -2860 362 -2855
rect 367 -2859 640 -2855
rect 367 -2860 571 -2859
rect 667 -2863 671 -2853
rect 659 -2909 663 -2903
rect 684 -2909 689 -2853
rect 694 -2852 697 -2848
rect 701 -2852 714 -2848
rect 718 -2852 721 -2848
rect 694 -2854 721 -2852
rect 702 -2859 706 -2854
rect 710 -2909 714 -2899
rect 855 -2909 860 -2648
rect 902 -2649 971 -2648
rect 993 -2678 997 -2672
rect 1018 -2678 1023 -2622
rect 1028 -2621 1031 -2617
rect 1035 -2621 1048 -2617
rect 1052 -2621 1055 -2617
rect 1028 -2623 1055 -2621
rect 1036 -2628 1040 -2623
rect 1044 -2678 1048 -2668
rect 993 -2682 1007 -2678
rect 1001 -2683 1007 -2682
rect 1018 -2683 1036 -2678
rect 1044 -2683 1202 -2678
rect 659 -2913 673 -2909
rect 667 -2914 673 -2913
rect 684 -2914 702 -2909
rect 710 -2914 860 -2909
rect 892 -2694 993 -2689
rect 568 -2921 659 -2920
rect 343 -2926 344 -2921
rect 349 -2925 659 -2921
rect 349 -2926 571 -2925
rect 667 -2928 671 -2914
rect 710 -2917 714 -2914
rect 702 -2943 706 -2937
rect 694 -2944 721 -2943
rect 694 -2948 695 -2944
rect 699 -2948 716 -2944
rect 720 -2948 721 -2944
rect 694 -2949 721 -2948
rect 659 -2974 663 -2968
rect 651 -2975 678 -2974
rect 651 -2979 652 -2975
rect 656 -2979 673 -2975
rect 677 -2979 678 -2975
rect 651 -2980 678 -2979
rect 892 -2994 897 -2694
rect 1001 -2697 1005 -2683
rect 1044 -2686 1048 -2683
rect 1036 -2712 1040 -2706
rect 1028 -2713 1055 -2712
rect 1028 -2717 1029 -2713
rect 1033 -2717 1050 -2713
rect 1054 -2717 1055 -2713
rect 1028 -2718 1055 -2717
rect 993 -2743 997 -2737
rect 985 -2744 1012 -2743
rect 985 -2748 986 -2744
rect 990 -2748 1007 -2744
rect 1011 -2748 1012 -2744
rect 985 -2749 1012 -2748
rect 967 -2830 1021 -2827
rect 967 -2834 970 -2830
rect 974 -2834 987 -2830
rect 991 -2834 997 -2830
rect 1001 -2834 1014 -2830
rect 1018 -2834 1021 -2830
rect 967 -2836 1021 -2834
rect 975 -2841 979 -2836
rect 1002 -2841 1006 -2836
rect 983 -2901 987 -2881
rect 1010 -2901 1014 -2881
rect 1029 -2900 1056 -2897
rect 983 -2905 1024 -2901
rect 568 -2995 897 -2994
rect 334 -3000 335 -2995
rect 340 -2999 897 -2995
rect 903 -2911 975 -2906
rect 340 -3000 571 -2999
rect 903 -3012 908 -2911
rect 1002 -2915 1006 -2905
rect 994 -2961 998 -2955
rect 1019 -2961 1024 -2905
rect 1029 -2904 1032 -2900
rect 1036 -2904 1049 -2900
rect 1053 -2904 1056 -2900
rect 1029 -2906 1056 -2904
rect 1037 -2911 1041 -2906
rect 1045 -2961 1049 -2951
rect 994 -2965 1008 -2961
rect 1002 -2966 1008 -2965
rect 1019 -2966 1037 -2961
rect 1045 -2966 1185 -2961
rect 736 -3017 908 -3012
rect 920 -2977 994 -2972
rect 628 -3049 682 -3046
rect 628 -3053 631 -3049
rect 635 -3053 648 -3049
rect 652 -3053 658 -3049
rect 662 -3053 675 -3049
rect 679 -3053 682 -3049
rect 628 -3055 682 -3053
rect 636 -3060 640 -3055
rect 663 -3060 667 -3055
rect 644 -3120 648 -3100
rect 671 -3120 675 -3100
rect 690 -3119 717 -3116
rect 644 -3124 685 -3120
rect 568 -3126 636 -3125
rect 367 -3130 636 -3126
rect 367 -3131 571 -3130
rect 663 -3134 667 -3124
rect 655 -3180 659 -3174
rect 680 -3180 685 -3124
rect 690 -3123 693 -3119
rect 697 -3123 710 -3119
rect 714 -3123 717 -3119
rect 690 -3125 717 -3123
rect 698 -3130 702 -3125
rect 706 -3180 710 -3170
rect 736 -3180 741 -3017
rect 920 -3034 925 -2977
rect 1002 -2980 1006 -2966
rect 1045 -2969 1049 -2966
rect 1037 -2995 1041 -2989
rect 1029 -2996 1056 -2995
rect 1029 -3000 1030 -2996
rect 1034 -3000 1051 -2996
rect 1055 -3000 1056 -2996
rect 1029 -3001 1056 -3000
rect 994 -3026 998 -3020
rect 986 -3027 1013 -3026
rect 986 -3031 987 -3027
rect 991 -3031 1008 -3027
rect 1012 -3031 1013 -3027
rect 986 -3032 1013 -3031
rect 655 -3184 669 -3180
rect 663 -3185 669 -3184
rect 680 -3185 698 -3180
rect 706 -3185 741 -3180
rect 750 -3039 925 -3034
rect 568 -3192 655 -3191
rect 343 -3197 344 -3192
rect 349 -3196 655 -3192
rect 349 -3197 571 -3196
rect 663 -3199 667 -3185
rect 706 -3188 710 -3185
rect 698 -3214 702 -3208
rect 690 -3215 717 -3214
rect 690 -3219 691 -3215
rect 695 -3219 712 -3215
rect 716 -3219 717 -3215
rect 690 -3220 717 -3219
rect 655 -3245 659 -3239
rect 647 -3246 674 -3245
rect 647 -3250 648 -3246
rect 652 -3250 669 -3246
rect 673 -3250 674 -3246
rect 647 -3251 674 -3250
rect 616 -3298 670 -3295
rect 616 -3302 619 -3298
rect 623 -3302 636 -3298
rect 640 -3302 646 -3298
rect 650 -3302 663 -3298
rect 667 -3302 670 -3298
rect 616 -3304 670 -3302
rect 624 -3309 628 -3304
rect 651 -3309 655 -3304
rect 632 -3369 636 -3349
rect 659 -3369 663 -3349
rect 678 -3368 705 -3365
rect 632 -3373 673 -3369
rect 568 -3375 624 -3374
rect 322 -3379 624 -3375
rect 322 -3380 571 -3379
rect 651 -3383 655 -3373
rect 643 -3429 647 -3423
rect 668 -3429 673 -3373
rect 678 -3372 681 -3368
rect 685 -3372 698 -3368
rect 702 -3372 705 -3368
rect 678 -3374 705 -3372
rect 686 -3379 690 -3374
rect 694 -3429 698 -3419
rect 750 -3429 755 -3039
rect 1180 -3074 1185 -2966
rect 1197 -2971 1202 -2683
rect 1213 -2685 1218 -2490
rect 1243 -2582 1248 -2459
rect 1296 -2488 1323 -2485
rect 1296 -2492 1299 -2488
rect 1303 -2492 1316 -2488
rect 1320 -2492 1323 -2488
rect 1296 -2494 1323 -2492
rect 1304 -2499 1308 -2494
rect 1243 -2587 1304 -2582
rect 1243 -2588 1248 -2587
rect 1312 -2591 1316 -2579
rect 1304 -2595 1316 -2591
rect 1304 -2599 1308 -2595
rect 1345 -2625 1372 -2622
rect 1345 -2629 1348 -2625
rect 1352 -2629 1365 -2625
rect 1369 -2629 1372 -2625
rect 1345 -2631 1372 -2629
rect 1353 -2636 1357 -2631
rect 1213 -2690 1289 -2685
rect 1312 -2686 1316 -2679
rect 1361 -2686 1365 -2676
rect 1312 -2691 1353 -2686
rect 1361 -2691 1445 -2686
rect 1312 -2694 1316 -2691
rect 1361 -2694 1365 -2691
rect 1297 -2698 1334 -2694
rect 1297 -2704 1301 -2698
rect 1330 -2704 1334 -2698
rect 1353 -2720 1357 -2714
rect 1345 -2721 1372 -2720
rect 1289 -2730 1293 -2724
rect 1322 -2730 1326 -2724
rect 1345 -2725 1346 -2721
rect 1350 -2725 1367 -2721
rect 1371 -2725 1372 -2721
rect 1345 -2726 1372 -2725
rect 1281 -2731 1308 -2730
rect 1281 -2735 1282 -2731
rect 1286 -2735 1303 -2731
rect 1307 -2735 1308 -2731
rect 1281 -2736 1308 -2735
rect 1314 -2731 1341 -2730
rect 1314 -2735 1315 -2731
rect 1319 -2735 1336 -2731
rect 1340 -2735 1341 -2731
rect 1314 -2736 1341 -2735
rect 1303 -2877 1330 -2874
rect 1303 -2881 1306 -2877
rect 1310 -2881 1323 -2877
rect 1327 -2881 1330 -2877
rect 1303 -2883 1330 -2881
rect 1311 -2888 1315 -2883
rect 1437 -2894 1445 -2691
rect 1800 -2802 1827 -2799
rect 1800 -2806 1803 -2802
rect 1807 -2806 1820 -2802
rect 1824 -2806 1827 -2802
rect 1800 -2808 1827 -2806
rect 1808 -2813 1812 -2808
rect 2272 -2828 2336 -2825
rect 2272 -2832 2275 -2828
rect 2279 -2832 2297 -2828
rect 2301 -2832 2307 -2828
rect 2311 -2832 2329 -2828
rect 2333 -2832 2336 -2828
rect 2071 -2836 2259 -2833
rect 2272 -2834 2336 -2832
rect 2071 -2840 2074 -2836
rect 2078 -2840 2096 -2836
rect 2100 -2840 2126 -2836
rect 2130 -2840 2148 -2836
rect 2152 -2840 2178 -2836
rect 2182 -2840 2200 -2836
rect 2204 -2840 2230 -2836
rect 2234 -2840 2252 -2836
rect 2256 -2840 2259 -2836
rect 2071 -2842 2259 -2840
rect 2282 -2840 2286 -2834
rect 2314 -2840 2318 -2834
rect 2081 -2848 2085 -2842
rect 2133 -2848 2137 -2842
rect 2185 -2848 2189 -2842
rect 2237 -2848 2241 -2842
rect 1437 -2897 1752 -2894
rect 1791 -2897 1808 -2896
rect 1437 -2901 1808 -2897
rect 1437 -2902 1793 -2901
rect 1437 -2904 1752 -2902
rect 1437 -2905 1730 -2904
rect 1816 -2905 1820 -2893
rect 1197 -2976 1311 -2971
rect 1319 -2980 1323 -2968
rect 1311 -2984 1323 -2980
rect 1808 -2909 1820 -2905
rect 2058 -2897 2081 -2892
rect 1808 -2913 1812 -2909
rect 2058 -2912 2063 -2897
rect 2089 -2901 2093 -2888
rect 1311 -2988 1315 -2984
rect 2032 -2920 2063 -2912
rect 1849 -2939 1876 -2936
rect 1849 -2943 1852 -2939
rect 1856 -2943 1869 -2939
rect 1873 -2943 1876 -2939
rect 1849 -2945 1876 -2943
rect 1857 -2950 1861 -2945
rect 1684 -2997 1692 -2996
rect 1684 -3000 1740 -2997
rect 1784 -3000 1793 -2999
rect 1684 -3004 1793 -3000
rect 1816 -3000 1820 -2993
rect 1865 -3000 1869 -2990
rect 2032 -2997 2039 -2920
rect 2058 -2963 2063 -2920
rect 2081 -2905 2093 -2901
rect 2111 -2897 2133 -2892
rect 2081 -2910 2085 -2905
rect 2076 -2959 2081 -2954
rect 2089 -2963 2093 -2950
rect 2111 -2963 2116 -2897
rect 2141 -2901 2145 -2888
rect 2193 -2892 2197 -2888
rect 2245 -2892 2249 -2888
rect 2290 -2892 2294 -2880
rect 2322 -2892 2326 -2880
rect 2133 -2905 2145 -2901
rect 2163 -2897 2185 -2892
rect 2193 -2897 2237 -2892
rect 2245 -2897 2282 -2892
rect 2290 -2897 2314 -2892
rect 2322 -2897 2336 -2892
rect 2133 -2910 2137 -2905
rect 2128 -2959 2133 -2954
rect 2141 -2963 2145 -2950
rect 2163 -2963 2168 -2897
rect 2182 -2920 2185 -2915
rect 2193 -2924 2197 -2897
rect 2185 -2955 2189 -2944
rect 2185 -2959 2197 -2955
rect 2058 -2968 2081 -2963
rect 2089 -2968 2133 -2963
rect 2141 -2968 2185 -2963
rect 2089 -2971 2093 -2968
rect 2141 -2971 2145 -2968
rect 2193 -2971 2197 -2959
rect 2215 -2963 2220 -2897
rect 2234 -2920 2237 -2915
rect 2245 -2924 2249 -2897
rect 2290 -2900 2294 -2897
rect 2322 -2900 2326 -2897
rect 2282 -2927 2286 -2920
rect 2314 -2927 2318 -2920
rect 2272 -2929 2336 -2927
rect 2272 -2933 2274 -2929
rect 2278 -2933 2298 -2929
rect 2302 -2933 2306 -2929
rect 2310 -2933 2330 -2929
rect 2334 -2933 2336 -2929
rect 2272 -2935 2336 -2933
rect 2237 -2955 2241 -2944
rect 2237 -2959 2249 -2955
rect 2215 -2968 2237 -2963
rect 2245 -2971 2249 -2959
rect 1881 -3000 2040 -2997
rect 2081 -2999 2085 -2991
rect 2133 -2999 2137 -2991
rect 2185 -2999 2189 -2991
rect 2237 -2999 2241 -2991
rect 1684 -3005 1786 -3004
rect 1816 -3005 1857 -3000
rect 1865 -3005 2040 -3000
rect 2071 -3000 2259 -2999
rect 2071 -3004 2098 -3000
rect 2102 -3004 2150 -3000
rect 2154 -3004 2202 -3000
rect 2206 -3004 2254 -3000
rect 2258 -3004 2259 -3000
rect 2071 -3005 2259 -3004
rect 1352 -3014 1379 -3011
rect 1352 -3018 1355 -3014
rect 1359 -3018 1372 -3014
rect 1376 -3018 1379 -3014
rect 1352 -3020 1379 -3018
rect 1360 -3025 1364 -3020
rect 1595 -3033 1622 -3030
rect 1595 -3037 1598 -3033
rect 1602 -3037 1615 -3033
rect 1619 -3037 1622 -3033
rect 1595 -3039 1622 -3037
rect 1180 -3079 1296 -3074
rect 1319 -3075 1323 -3068
rect 1368 -3075 1372 -3065
rect 1603 -3044 1607 -3039
rect 1319 -3080 1360 -3075
rect 1368 -3080 1573 -3075
rect 1319 -3083 1323 -3080
rect 1368 -3083 1372 -3080
rect 1304 -3087 1341 -3083
rect 1304 -3093 1308 -3087
rect 1337 -3093 1341 -3087
rect 1360 -3109 1364 -3103
rect 1352 -3110 1379 -3109
rect 1296 -3119 1300 -3113
rect 1329 -3119 1333 -3113
rect 1352 -3114 1353 -3110
rect 1357 -3114 1374 -3110
rect 1378 -3114 1379 -3110
rect 1352 -3115 1379 -3114
rect 1288 -3120 1315 -3119
rect 1288 -3124 1289 -3120
rect 1293 -3124 1310 -3120
rect 1314 -3124 1315 -3120
rect 1288 -3125 1315 -3124
rect 1321 -3120 1348 -3119
rect 1321 -3124 1322 -3120
rect 1326 -3124 1343 -3120
rect 1347 -3124 1348 -3120
rect 1321 -3125 1348 -3124
rect 1568 -3128 1573 -3080
rect 1684 -3067 1692 -3005
rect 1816 -3008 1820 -3005
rect 1865 -3008 1869 -3005
rect 1801 -3012 1838 -3008
rect 1801 -3018 1805 -3012
rect 1834 -3018 1838 -3012
rect 2064 -3018 2071 -3013
rect 2076 -3018 2123 -3013
rect 2128 -3018 2177 -3013
rect 2182 -3018 2229 -3013
rect 1857 -3034 1861 -3028
rect 1849 -3035 1876 -3034
rect 1793 -3044 1797 -3038
rect 1826 -3044 1830 -3038
rect 1849 -3039 1850 -3035
rect 1854 -3039 1871 -3035
rect 1875 -3039 1876 -3035
rect 1849 -3040 1876 -3039
rect 1785 -3045 1812 -3044
rect 1785 -3049 1786 -3045
rect 1790 -3049 1807 -3045
rect 1811 -3049 1812 -3045
rect 1785 -3050 1812 -3049
rect 1818 -3045 1845 -3044
rect 1818 -3049 1819 -3045
rect 1823 -3049 1840 -3045
rect 1844 -3049 1845 -3045
rect 1818 -3050 1845 -3049
rect 1586 -3128 1603 -3127
rect 1568 -3132 1603 -3128
rect 1568 -3133 1592 -3132
rect 1611 -3136 1615 -3124
rect 1603 -3140 1615 -3136
rect 1603 -3144 1607 -3140
rect 1683 -3165 1692 -3067
rect 1644 -3170 1671 -3167
rect 1644 -3174 1647 -3170
rect 1651 -3174 1664 -3170
rect 1668 -3174 1671 -3170
rect 1644 -3176 1671 -3174
rect 1652 -3181 1656 -3176
rect 1297 -3232 1351 -3229
rect 1297 -3236 1300 -3232
rect 1304 -3236 1317 -3232
rect 1321 -3236 1327 -3232
rect 1331 -3236 1344 -3232
rect 1348 -3236 1351 -3232
rect 1297 -3238 1351 -3236
rect 1554 -3235 1588 -3230
rect 1611 -3231 1615 -3224
rect 1660 -3231 1664 -3221
rect 1683 -3231 1691 -3165
rect 1305 -3243 1309 -3238
rect 1332 -3243 1336 -3238
rect 1313 -3303 1317 -3283
rect 1340 -3303 1344 -3283
rect 1359 -3302 1386 -3299
rect 643 -3433 657 -3429
rect 651 -3434 657 -3433
rect 668 -3434 686 -3429
rect 694 -3434 755 -3429
rect 760 -3308 1302 -3304
rect 1313 -3307 1354 -3303
rect 760 -3309 1305 -3308
rect 568 -3441 643 -3440
rect 325 -3446 326 -3441
rect 331 -3445 643 -3441
rect 331 -3446 571 -3445
rect 651 -3448 655 -3434
rect 694 -3437 698 -3434
rect 686 -3463 690 -3457
rect 678 -3464 705 -3463
rect 678 -3468 679 -3464
rect 683 -3468 700 -3464
rect 704 -3468 705 -3464
rect 678 -3469 705 -3468
rect 643 -3494 647 -3488
rect 635 -3495 662 -3494
rect 635 -3499 636 -3495
rect 640 -3499 657 -3495
rect 661 -3499 662 -3495
rect 635 -3500 662 -3499
rect 633 -3565 687 -3562
rect 633 -3569 636 -3565
rect 640 -3569 653 -3565
rect 657 -3569 663 -3565
rect 667 -3569 680 -3565
rect 684 -3569 687 -3565
rect 633 -3571 687 -3569
rect 641 -3576 645 -3571
rect 668 -3576 672 -3571
rect 649 -3636 653 -3616
rect 676 -3636 680 -3616
rect 695 -3635 722 -3632
rect 649 -3640 690 -3636
rect 568 -3642 641 -3641
rect 298 -3647 299 -3642
rect 304 -3646 641 -3642
rect 304 -3647 571 -3646
rect 668 -3650 672 -3640
rect 660 -3696 664 -3690
rect 685 -3696 690 -3640
rect 695 -3639 698 -3635
rect 702 -3639 715 -3635
rect 719 -3639 722 -3635
rect 695 -3641 722 -3639
rect 703 -3646 707 -3641
rect 711 -3696 715 -3686
rect 760 -3696 765 -3309
rect 1297 -3313 1305 -3309
rect 1297 -3314 1302 -3313
rect 1332 -3317 1336 -3307
rect 957 -3364 1011 -3361
rect 957 -3368 960 -3364
rect 964 -3368 977 -3364
rect 981 -3368 987 -3364
rect 991 -3368 1004 -3364
rect 1008 -3368 1011 -3364
rect 1324 -3363 1328 -3357
rect 1349 -3363 1354 -3307
rect 1359 -3306 1362 -3302
rect 1366 -3306 1379 -3302
rect 1383 -3306 1386 -3302
rect 1359 -3308 1386 -3306
rect 1367 -3313 1371 -3308
rect 1375 -3363 1379 -3353
rect 1554 -3363 1559 -3235
rect 1611 -3236 1652 -3231
rect 1660 -3236 1691 -3231
rect 1611 -3239 1615 -3236
rect 1660 -3239 1664 -3236
rect 1596 -3243 1633 -3239
rect 1596 -3249 1600 -3243
rect 1629 -3249 1633 -3243
rect 1652 -3265 1656 -3259
rect 1644 -3266 1671 -3265
rect 1588 -3275 1592 -3269
rect 1621 -3275 1625 -3269
rect 1644 -3270 1645 -3266
rect 1649 -3270 1666 -3266
rect 1670 -3270 1671 -3266
rect 1644 -3271 1671 -3270
rect 1580 -3276 1607 -3275
rect 1580 -3280 1581 -3276
rect 1585 -3280 1602 -3276
rect 1606 -3280 1607 -3276
rect 1580 -3281 1607 -3280
rect 1613 -3276 1640 -3275
rect 1613 -3280 1614 -3276
rect 1618 -3280 1635 -3276
rect 1639 -3280 1640 -3276
rect 1613 -3281 1640 -3280
rect 1324 -3367 1338 -3363
rect 957 -3370 1011 -3368
rect 1332 -3368 1338 -3367
rect 1349 -3368 1367 -3363
rect 1375 -3368 1559 -3363
rect 965 -3375 969 -3370
rect 992 -3375 996 -3370
rect 973 -3435 977 -3415
rect 1000 -3435 1004 -3415
rect 1100 -3379 1324 -3374
rect 1019 -3434 1046 -3431
rect 958 -3440 963 -3438
rect 973 -3439 1014 -3435
rect 958 -3442 965 -3440
rect 660 -3700 674 -3696
rect 668 -3701 674 -3700
rect 685 -3701 703 -3696
rect 711 -3701 765 -3696
rect 845 -3445 965 -3442
rect 845 -3447 963 -3445
rect 568 -3708 660 -3707
rect 307 -3713 308 -3708
rect 313 -3712 660 -3708
rect 313 -3713 571 -3712
rect 668 -3715 672 -3701
rect 711 -3704 715 -3701
rect 703 -3730 707 -3724
rect 695 -3731 722 -3730
rect 695 -3735 696 -3731
rect 700 -3735 717 -3731
rect 721 -3735 722 -3731
rect 695 -3736 722 -3735
rect 660 -3761 664 -3755
rect 652 -3762 679 -3761
rect 652 -3766 653 -3762
rect 657 -3766 674 -3762
rect 678 -3766 679 -3762
rect 652 -3767 679 -3766
rect 621 -3814 675 -3811
rect 621 -3818 624 -3814
rect 628 -3818 641 -3814
rect 645 -3818 651 -3814
rect 655 -3818 668 -3814
rect 672 -3818 675 -3814
rect 621 -3820 675 -3818
rect 629 -3825 633 -3820
rect 656 -3825 660 -3820
rect 637 -3885 641 -3865
rect 664 -3885 668 -3865
rect 683 -3884 710 -3881
rect 637 -3889 678 -3885
rect 568 -3891 629 -3890
rect 325 -3896 326 -3891
rect 331 -3895 629 -3891
rect 331 -3896 571 -3895
rect 656 -3899 660 -3889
rect 648 -3945 652 -3939
rect 673 -3945 678 -3889
rect 683 -3888 686 -3884
rect 690 -3888 703 -3884
rect 707 -3888 710 -3884
rect 683 -3890 710 -3888
rect 691 -3895 695 -3890
rect 699 -3945 703 -3935
rect 845 -3945 850 -3447
rect 958 -3449 963 -3447
rect 992 -3449 996 -3439
rect 984 -3495 988 -3489
rect 1009 -3495 1014 -3439
rect 1019 -3438 1022 -3434
rect 1026 -3438 1039 -3434
rect 1043 -3438 1046 -3434
rect 1019 -3440 1046 -3438
rect 1027 -3445 1031 -3440
rect 1035 -3495 1039 -3485
rect 1100 -3494 1105 -3379
rect 1332 -3382 1336 -3368
rect 1375 -3371 1379 -3368
rect 1367 -3397 1371 -3391
rect 1359 -3398 1386 -3397
rect 1359 -3402 1360 -3398
rect 1364 -3402 1381 -3398
rect 1385 -3402 1386 -3398
rect 1359 -3403 1386 -3402
rect 1324 -3428 1328 -3422
rect 1316 -3429 1343 -3428
rect 1316 -3433 1317 -3429
rect 1321 -3433 1338 -3429
rect 1342 -3433 1343 -3429
rect 1316 -3434 1343 -3433
rect 1045 -3495 1105 -3494
rect 984 -3499 998 -3495
rect 992 -3500 998 -3499
rect 1009 -3500 1027 -3495
rect 1035 -3499 1105 -3495
rect 1035 -3500 1048 -3499
rect 648 -3949 662 -3945
rect 656 -3950 662 -3949
rect 673 -3950 691 -3945
rect 699 -3950 850 -3945
rect 891 -3511 984 -3506
rect 568 -3957 648 -3956
rect 343 -3962 344 -3957
rect 349 -3961 648 -3957
rect 349 -3962 571 -3961
rect 656 -3964 660 -3950
rect 699 -3953 703 -3950
rect 691 -3979 695 -3973
rect 683 -3980 710 -3979
rect 683 -3984 684 -3980
rect 688 -3984 705 -3980
rect 709 -3984 710 -3980
rect 683 -3985 710 -3984
rect 648 -4010 652 -4004
rect 640 -4011 667 -4010
rect 640 -4015 641 -4011
rect 645 -4015 662 -4011
rect 666 -4015 667 -4011
rect 640 -4016 667 -4015
rect 891 -4025 896 -3511
rect 992 -3514 996 -3500
rect 1035 -3503 1039 -3500
rect 1027 -3529 1031 -3523
rect 1019 -3530 1046 -3529
rect 1019 -3534 1020 -3530
rect 1024 -3534 1041 -3530
rect 1045 -3534 1046 -3530
rect 1019 -3535 1046 -3534
rect 984 -3560 988 -3554
rect 976 -3561 1003 -3560
rect 976 -3565 977 -3561
rect 981 -3565 998 -3561
rect 1002 -3565 1003 -3561
rect 976 -3566 1003 -3565
rect 568 -4026 896 -4025
rect 361 -4031 362 -4026
rect 367 -4030 896 -4026
rect 367 -4031 571 -4030
<< m2contact >>
rect -1538 288 -1533 293
rect -1486 288 -1481 293
rect -1432 327 -1427 332
rect -1380 327 -1375 332
rect 3757 285 3762 290
rect 3809 285 3814 290
rect 3863 324 3868 329
rect 3915 324 3920 329
rect -1538 229 -1533 234
rect -1486 229 -1481 234
rect -1432 229 -1427 234
rect -1380 229 -1375 234
rect 3757 226 3762 231
rect 3809 226 3814 231
rect 3863 226 3868 231
rect 3915 226 3920 231
rect 299 26 304 31
rect 308 -22 313 -17
rect 1409 -18 1414 -13
rect -412 -113 -407 -108
rect -360 -113 -355 -108
rect -306 -74 -301 -69
rect -254 -74 -249 -69
rect -412 -172 -407 -167
rect -360 -172 -355 -167
rect -306 -172 -301 -167
rect -254 -172 -249 -167
rect 1461 -18 1466 -13
rect 1515 21 1520 26
rect 1567 21 1572 26
rect 1409 -77 1414 -72
rect 1461 -77 1466 -72
rect 1515 -77 1520 -72
rect 1567 -77 1572 -72
rect 14 -176 19 -171
rect 308 -218 313 -213
rect -416 -368 -411 -363
rect -364 -368 -359 -363
rect -310 -329 -305 -324
rect -258 -329 -253 -324
rect -416 -427 -411 -422
rect -364 -427 -359 -422
rect -310 -427 -305 -422
rect -258 -427 -253 -422
rect 299 -284 304 -279
rect 101 -377 107 -372
rect 317 -432 322 -427
rect 326 -461 331 -456
rect 1424 -294 1429 -289
rect 1476 -294 1481 -289
rect 1530 -255 1535 -250
rect 1582 -255 1587 -250
rect 1424 -353 1429 -348
rect 1476 -353 1481 -348
rect 1530 -353 1535 -348
rect 1582 -353 1587 -348
rect 335 -864 340 -859
rect -319 -950 -314 -945
rect 317 -888 322 -883
rect -267 -950 -262 -945
rect -213 -911 -208 -906
rect -161 -911 -156 -906
rect 2 -962 7 -957
rect -319 -1009 -314 -1004
rect -267 -1009 -262 -1004
rect -213 -1009 -208 -1004
rect -161 -1009 -156 -1004
rect 326 -1004 331 -999
rect -338 -1173 -333 -1168
rect -286 -1173 -281 -1168
rect -232 -1134 -227 -1129
rect -180 -1134 -175 -1129
rect 299 -1133 304 -1128
rect 308 -1145 313 -1140
rect 89 -1163 95 -1158
rect 335 -1218 340 -1213
rect -338 -1232 -333 -1227
rect -286 -1232 -281 -1227
rect -232 -1232 -227 -1227
rect -180 -1232 -175 -1227
rect 1808 -967 1813 -962
rect 1860 -967 1865 -962
rect 1914 -928 1919 -923
rect 1966 -928 1971 -923
rect 1808 -1026 1813 -1021
rect 1860 -1026 1865 -1021
rect 1914 -1026 1919 -1021
rect 1966 -1026 1971 -1021
rect 326 -1271 331 -1266
rect 344 -1305 349 -1299
rect 353 -1319 358 -1314
rect 344 -1425 349 -1420
rect -338 -1511 -333 -1506
rect -286 -1511 -281 -1506
rect -232 -1472 -227 -1467
rect -180 -1472 -175 -1467
rect -338 -1570 -333 -1565
rect -286 -1570 -281 -1565
rect -232 -1570 -227 -1565
rect -180 -1570 -175 -1565
rect 335 -1491 340 -1486
rect 11 -1622 16 -1617
rect 344 -1664 349 -1659
rect -353 -1848 -348 -1843
rect -301 -1848 -296 -1843
rect -247 -1809 -242 -1804
rect -195 -1809 -190 -1804
rect 344 -1708 349 -1703
rect 326 -1774 331 -1769
rect 98 -1823 104 -1818
rect 317 -1845 322 -1840
rect 353 -1878 358 -1873
rect -353 -1907 -348 -1902
rect -301 -1907 -296 -1902
rect -247 -1907 -242 -1902
rect -195 -1907 -190 -1902
rect 299 -1979 304 -1974
rect 308 -2045 313 -2040
rect 1997 -1717 2002 -1712
rect 2049 -1717 2054 -1712
rect 2103 -1678 2108 -1673
rect 2155 -1678 2160 -1673
rect 1997 -1776 2002 -1771
rect 2049 -1776 2054 -1771
rect 2103 -1776 2108 -1771
rect 2155 -1776 2160 -1771
rect 344 -2228 349 -2223
rect 326 -2294 331 -2289
rect -353 -2455 -348 -2450
rect 362 -2383 367 -2378
rect -301 -2455 -296 -2450
rect -247 -2416 -242 -2411
rect -195 -2416 -190 -2411
rect 8 -2497 13 -2492
rect -353 -2514 -348 -2509
rect -301 -2514 -296 -2509
rect -247 -2514 -242 -2509
rect -195 -2514 -190 -2509
rect 362 -2539 367 -2534
rect -353 -2725 -348 -2720
rect -301 -2725 -296 -2720
rect -247 -2686 -242 -2681
rect -195 -2686 -190 -2681
rect 95 -2698 101 -2693
rect -353 -2784 -348 -2779
rect -301 -2784 -296 -2779
rect -247 -2784 -242 -2779
rect -195 -2784 -190 -2779
rect 353 -2770 358 -2765
rect 362 -2779 367 -2774
rect 362 -2860 367 -2855
rect 344 -2926 349 -2921
rect 335 -3000 340 -2995
rect 362 -3131 367 -3126
rect 344 -3197 349 -3192
rect 317 -3380 322 -3375
rect 2071 -2959 2076 -2954
rect 2123 -2959 2128 -2954
rect 2177 -2920 2182 -2915
rect 2229 -2920 2234 -2915
rect 2071 -3018 2076 -3013
rect 2123 -3018 2128 -3013
rect 2177 -3018 2182 -3013
rect 2229 -3018 2234 -3013
rect 326 -3446 331 -3441
rect 299 -3647 304 -3642
rect 308 -3713 313 -3708
rect 326 -3896 331 -3891
rect 344 -3962 349 -3957
rect 362 -4031 367 -4026
<< metal2 >>
rect -1538 234 -1533 288
rect -1486 234 -1481 288
rect -1432 234 -1427 327
rect -1380 234 -1375 327
rect 3757 231 3762 285
rect 3809 231 3814 285
rect 3863 231 3868 324
rect 3915 231 3920 324
rect -412 -167 -407 -113
rect -360 -167 -355 -113
rect -306 -167 -301 -74
rect -254 -167 -249 -74
rect -416 -422 -411 -368
rect -364 -422 -359 -368
rect -310 -422 -305 -329
rect -258 -422 -253 -329
rect 14 -372 19 -176
rect 299 -279 304 26
rect 14 -377 101 -372
rect -319 -1004 -314 -950
rect -267 -1004 -262 -950
rect -213 -1004 -208 -911
rect -161 -1004 -156 -911
rect -338 -1227 -333 -1173
rect -286 -1227 -281 -1173
rect -232 -1227 -227 -1134
rect -180 -1227 -175 -1134
rect 2 -1158 7 -962
rect 299 -1128 304 -284
rect 2 -1163 89 -1158
rect -338 -1565 -333 -1511
rect -286 -1565 -281 -1511
rect -232 -1565 -227 -1472
rect -180 -1565 -175 -1472
rect -353 -1902 -348 -1848
rect -301 -1902 -296 -1848
rect -247 -1902 -242 -1809
rect -195 -1902 -190 -1809
rect 11 -1818 16 -1622
rect 11 -1823 98 -1818
rect 299 -1974 304 -1133
rect -353 -2509 -348 -2455
rect -301 -2509 -296 -2455
rect -247 -2509 -242 -2416
rect -195 -2509 -190 -2416
rect -353 -2779 -348 -2725
rect -301 -2779 -296 -2725
rect -247 -2779 -242 -2686
rect -195 -2779 -190 -2686
rect 8 -2693 13 -2497
rect 8 -2698 95 -2693
rect 299 -3642 304 -1979
rect 299 -4035 304 -3647
rect 308 -213 313 -22
rect 1409 -72 1414 -18
rect 1461 -72 1466 -18
rect 1515 -72 1520 21
rect 1567 -72 1572 21
rect 308 -1140 313 -218
rect 1424 -348 1429 -294
rect 1476 -348 1481 -294
rect 1530 -348 1535 -255
rect 1582 -348 1587 -255
rect 308 -2040 313 -1145
rect 308 -3708 313 -2045
rect 308 -4036 313 -3713
rect 317 -883 322 -432
rect 317 -1840 322 -888
rect 317 -3375 322 -1845
rect 317 -4032 322 -3380
rect 326 -999 331 -461
rect 326 -1266 331 -1004
rect 326 -1769 331 -1271
rect 326 -2289 331 -1774
rect 326 -3441 331 -2294
rect 326 -3891 331 -3446
rect 326 -4034 331 -3896
rect 335 -1213 340 -864
rect 1808 -1021 1813 -967
rect 1860 -1021 1865 -967
rect 1914 -1021 1919 -928
rect 1966 -1021 1971 -928
rect 335 -1486 340 -1218
rect 335 -2995 340 -1491
rect 335 -4033 340 -3000
rect 344 -1420 349 -1305
rect 344 -1659 349 -1425
rect 344 -1703 349 -1664
rect 344 -2223 349 -1708
rect 344 -2921 349 -2228
rect 344 -3192 349 -2926
rect 344 -3957 349 -3197
rect 344 -4033 349 -3962
rect 353 -1873 358 -1319
rect 1997 -1771 2002 -1717
rect 2049 -1771 2054 -1717
rect 2103 -1771 2108 -1678
rect 2155 -1771 2160 -1678
rect 353 -2765 358 -1878
rect 353 -4034 358 -2770
rect 362 -2378 367 -2373
rect 362 -2534 367 -2383
rect 362 -2774 367 -2539
rect 362 -2855 367 -2779
rect 362 -3126 367 -2860
rect 2071 -3013 2076 -2959
rect 2123 -3013 2128 -2959
rect 2177 -3013 2182 -2920
rect 2229 -3013 2234 -2920
rect 362 -4026 367 -3131
rect 362 -4034 367 -4031
<< labels >>
rlabel metal1 207 -243 207 -243 7 vdd
rlabel metal1 111 -243 111 -243 3 gnd
rlabel metal1 207 -192 207 -192 7 vdd
rlabel metal1 111 -192 111 -192 3 gnd
rlabel metal1 259 -250 259 -250 1 gnd
rlabel metal1 259 -154 259 -154 5 vdd
rlabel metal1 176 -298 176 -298 5 vdd
rlabel metal1 203 -298 203 -298 5 vdd
rlabel metal1 195 -495 195 -495 1 gnd
rlabel metal1 238 -368 238 -368 5 vdd
rlabel metal1 238 -464 238 -464 1 gnd
rlabel metal1 292 -430 292 -430 1 G0
rlabel metal1 287 -216 287 -216 1 P0
rlabel metal1 204 -1689 204 -1689 7 vdd
rlabel metal1 108 -1689 108 -1689 3 gnd
rlabel metal1 204 -1638 204 -1638 7 vdd
rlabel metal1 108 -1638 108 -1638 3 gnd
rlabel metal1 256 -1696 256 -1696 1 gnd
rlabel metal1 256 -1600 256 -1600 5 vdd
rlabel metal1 173 -1744 173 -1744 5 vdd
rlabel metal1 200 -1744 200 -1744 5 vdd
rlabel metal1 192 -1941 192 -1941 1 gnd
rlabel metal1 235 -1814 235 -1814 5 vdd
rlabel metal1 235 -1910 235 -1910 1 gnd
rlabel metal1 290 -1662 290 -1662 1 P2
rlabel metal1 287 -1876 287 -1876 1 G2
rlabel metal1 195 -1029 195 -1029 7 vdd
rlabel metal1 99 -1029 99 -1029 3 gnd
rlabel metal1 195 -978 195 -978 7 vdd
rlabel metal1 99 -978 99 -978 3 gnd
rlabel metal1 247 -1036 247 -1036 1 gnd
rlabel metal1 247 -940 247 -940 5 vdd
rlabel metal1 164 -1084 164 -1084 5 vdd
rlabel metal1 191 -1084 191 -1084 5 vdd
rlabel metal1 183 -1281 183 -1281 1 gnd
rlabel metal1 226 -1154 226 -1154 5 vdd
rlabel metal1 226 -1250 226 -1250 1 gnd
rlabel metal1 281 -1002 281 -1002 1 P1
rlabel metal1 281 -1216 281 -1216 1 G1
rlabel metal1 201 -2564 201 -2564 7 vdd
rlabel metal1 105 -2564 105 -2564 3 gnd
rlabel metal1 201 -2513 201 -2513 7 vdd
rlabel metal1 105 -2513 105 -2513 3 gnd
rlabel metal1 253 -2571 253 -2571 1 gnd
rlabel metal1 253 -2475 253 -2475 5 vdd
rlabel metal1 170 -2619 170 -2619 5 vdd
rlabel metal1 197 -2619 197 -2619 5 vdd
rlabel metal1 189 -2816 189 -2816 1 gnd
rlabel metal1 232 -2689 232 -2689 5 vdd
rlabel metal1 232 -2785 232 -2785 1 gnd
rlabel metal1 287 -2537 287 -2537 1 P3
rlabel metal1 284 -2751 284 -2751 1 G3
rlabel metal1 -14 28 -14 28 1 c0
rlabel metal1 -3492 -1263 -3492 -1263 7 vdd
rlabel metal1 -3588 -1263 -3588 -1263 3 gnd
rlabel metal1 -3492 -1212 -3492 -1212 7 vdd
rlabel metal1 -3588 -1212 -3588 -1212 3 gnd
rlabel metal1 -3440 -1270 -3440 -1270 1 gnd
rlabel metal1 -3440 -1174 -3440 -1174 5 vdd
rlabel metal1 -3113 -1325 -3113 -1325 1 gnd
rlabel metal1 -3113 -1229 -3113 -1229 5 vdd
rlabel metal1 -3156 -1356 -3156 -1356 1 gnd
rlabel metal1 -3148 -1159 -3148 -1159 5 vdd
rlabel metal1 -3175 -1159 -3175 -1159 5 vdd
rlabel metal1 -3235 -1380 -3235 -1380 1 gnd
rlabel metal1 -3235 -1284 -3235 -1284 5 vdd
rlabel metal1 -3266 -1390 -3266 -1390 1 gnd
rlabel metal1 -3299 -1390 -3299 -1390 1 gnd
rlabel metal1 -3284 -1147 -3284 -1147 5 vdd
rlabel metal1 -3349 -1286 -3349 -1286 1 gnd
rlabel metal1 -3349 -1190 -3349 -1190 5 vdd
rlabel metal1 821 -51 821 -51 5 vdd
rlabel metal1 806 -294 806 -294 1 gnd
rlabel metal1 839 -294 839 -294 1 gnd
rlabel metal1 870 -188 870 -188 5 vdd
rlabel metal1 870 -284 870 -284 1 gnd
rlabel metal1 513 -302 513 -302 1 gnd
rlabel metal1 513 -206 513 -206 5 vdd
rlabel metal1 470 -333 470 -333 1 gnd
rlabel metal1 478 -136 478 -136 5 vdd
rlabel metal1 451 -136 451 -136 5 vdd
rlabel metal1 890 -248 890 -248 1 c1
rlabel metal1 772 -1032 772 -1032 5 vdd
rlabel metal1 799 -1032 799 -1032 5 vdd
rlabel metal1 791 -1229 791 -1229 1 gnd
rlabel metal1 834 -1102 834 -1102 5 vdd
rlabel metal1 834 -1198 834 -1198 1 gnd
rlabel metal1 554 -1032 554 -1032 5 vdd
rlabel metal1 581 -1032 581 -1032 5 vdd
rlabel metal1 573 -1229 573 -1229 1 gnd
rlabel metal1 616 -1102 616 -1102 5 vdd
rlabel metal1 616 -1198 616 -1198 1 gnd
rlabel metal1 631 -787 631 -787 5 vdd
rlabel metal1 658 -787 658 -787 5 vdd
rlabel metal1 650 -984 650 -984 1 gnd
rlabel metal1 693 -857 693 -857 5 vdd
rlabel metal1 693 -953 693 -953 1 gnd
rlabel metal1 965 -698 965 -698 5 vdd
rlabel metal1 950 -941 950 -941 1 gnd
rlabel metal1 983 -941 983 -941 1 gnd
rlabel metal1 1014 -835 1014 -835 5 vdd
rlabel metal1 1014 -931 1014 -931 1 gnd
rlabel metal1 1216 -700 1216 -700 5 vdd
rlabel metal1 1201 -943 1201 -943 1 gnd
rlabel metal1 1234 -943 1234 -943 1 gnd
rlabel metal1 1265 -837 1265 -837 5 vdd
rlabel metal1 1265 -933 1265 -933 1 gnd
rlabel metal1 1619 -905 1619 -905 5 vdd
rlabel metal1 1619 -1001 1619 -1001 1 gnd
rlabel metal1 1471 -943 1471 -943 3 gnd
rlabel metal1 1567 -943 1567 -943 7 vdd
rlabel metal1 1471 -994 1471 -994 3 gnd
rlabel metal1 1567 -994 1567 -994 7 vdd
rlabel metal1 1167 -175 1167 -175 5 vdd
rlabel metal1 1167 -271 1167 -271 1 gnd
rlabel metal1 1019 -213 1019 -213 3 gnd
rlabel metal1 1115 -213 1115 -213 7 vdd
rlabel metal1 1019 -264 1019 -264 3 gnd
rlabel metal1 1115 -264 1115 -264 7 vdd
rlabel metal1 1172 45 1172 45 5 vdd
rlabel metal1 1172 -51 1172 -51 1 gnd
rlabel metal1 1024 7 1024 7 3 gnd
rlabel metal1 1120 7 1120 7 7 vdd
rlabel metal1 1024 -44 1024 -44 3 gnd
rlabel metal1 1120 -44 1120 -44 7 vdd
rlabel metal1 563 -1901 563 -1901 5 vdd
rlabel metal1 865 -1743 865 -1743 1 gnd
rlabel metal1 570 -2347 570 -2347 1 gnd
rlabel metal1 551 -2150 551 -2150 5 vdd
rlabel metal1 578 -2150 578 -2150 5 vdd
rlabel metal1 613 -2220 613 -2220 5 vdd
rlabel metal1 613 -2316 613 -2316 1 gnd
rlabel metal1 566 -1347 566 -1347 5 vdd
rlabel metal1 593 -1347 593 -1347 5 vdd
rlabel metal1 585 -1544 585 -1544 1 gnd
rlabel metal1 628 -1417 628 -1417 5 vdd
rlabel metal1 628 -1513 628 -1513 1 gnd
rlabel metal1 567 -1630 567 -1630 5 vdd
rlabel metal1 594 -1630 594 -1630 5 vdd
rlabel metal1 586 -1827 586 -1827 1 gnd
rlabel metal1 629 -1700 629 -1700 5 vdd
rlabel metal1 629 -1796 629 -1796 1 gnd
rlabel metal1 590 -1901 590 -1901 5 vdd
rlabel metal1 582 -2098 582 -2098 1 gnd
rlabel metal1 625 -1971 625 -1971 5 vdd
rlabel metal1 625 -2067 625 -2067 1 gnd
rlabel metal1 812 -1788 812 -1788 5 vdd
rlabel metal1 839 -1788 839 -1788 5 vdd
rlabel metal1 831 -1985 831 -1985 1 gnd
rlabel metal1 874 -1858 874 -1858 5 vdd
rlabel metal1 874 -1954 874 -1954 1 gnd
rlabel metal1 803 -1577 803 -1577 5 vdd
rlabel metal1 830 -1577 830 -1577 5 vdd
rlabel metal1 822 -1774 822 -1774 1 gnd
rlabel metal1 865 -1647 865 -1647 5 vdd
rlabel metal1 1096 -1723 1096 -1723 5 vdd
rlabel metal1 1081 -1966 1081 -1966 1 gnd
rlabel metal1 1114 -1966 1114 -1966 1 gnd
rlabel metal1 1145 -1860 1145 -1860 5 vdd
rlabel metal1 1145 -1956 1145 -1956 1 gnd
rlabel metal1 1085 -1423 1085 -1423 5 vdd
rlabel metal1 1070 -1666 1070 -1666 1 gnd
rlabel metal1 1103 -1666 1103 -1666 1 gnd
rlabel metal1 1134 -1560 1134 -1560 5 vdd
rlabel metal1 1134 -1656 1134 -1656 1 gnd
rlabel metal1 1382 -1576 1382 -1576 5 vdd
rlabel metal1 1367 -1819 1367 -1819 1 gnd
rlabel metal1 1400 -1819 1400 -1819 1 gnd
rlabel metal1 1431 -1713 1431 -1713 5 vdd
rlabel metal1 1431 -1809 1431 -1809 1 gnd
rlabel metal1 1800 -1641 1800 -1641 5 vdd
rlabel metal1 1800 -1737 1800 -1737 1 gnd
rlabel metal1 1652 -1679 1652 -1679 3 gnd
rlabel metal1 1748 -1679 1748 -1679 7 vdd
rlabel metal1 1652 -1730 1652 -1730 3 gnd
rlabel metal1 1748 -1730 1748 -1730 7 vdd
rlabel metal1 1358 -2723 1358 -2723 1 gnd
rlabel metal1 1358 -2627 1358 -2627 5 vdd
rlabel metal1 1327 -2733 1327 -2733 1 gnd
rlabel metal1 1294 -2733 1294 -2733 1 gnd
rlabel metal1 1309 -2490 1309 -2490 5 vdd
rlabel metal1 1365 -3112 1365 -3112 1 gnd
rlabel metal1 1365 -3016 1365 -3016 5 vdd
rlabel metal1 1334 -3122 1334 -3122 1 gnd
rlabel metal1 1301 -3122 1301 -3122 1 gnd
rlabel metal1 1316 -2879 1316 -2879 5 vdd
rlabel metal1 1657 -3268 1657 -3268 1 gnd
rlabel metal1 1657 -3172 1657 -3172 5 vdd
rlabel metal1 1626 -3278 1626 -3278 1 gnd
rlabel metal1 1593 -3278 1593 -3278 1 gnd
rlabel metal1 1608 -3035 1608 -3035 5 vdd
rlabel metal1 703 -3217 703 -3217 1 gnd
rlabel metal1 703 -3121 703 -3121 5 vdd
rlabel metal1 660 -3248 660 -3248 1 gnd
rlabel metal1 668 -3051 668 -3051 5 vdd
rlabel metal1 641 -3051 641 -3051 5 vdd
rlabel metal1 707 -2946 707 -2946 1 gnd
rlabel metal1 707 -2850 707 -2850 5 vdd
rlabel metal1 664 -2977 664 -2977 1 gnd
rlabel metal1 672 -2780 672 -2780 5 vdd
rlabel metal1 645 -2780 645 -2780 5 vdd
rlabel metal1 706 -2663 706 -2663 1 gnd
rlabel metal1 706 -2567 706 -2567 5 vdd
rlabel metal1 663 -2694 663 -2694 1 gnd
rlabel metal1 671 -2497 671 -2497 5 vdd
rlabel metal1 644 -2497 644 -2497 5 vdd
rlabel metal1 691 -3466 691 -3466 1 gnd
rlabel metal1 691 -3370 691 -3370 5 vdd
rlabel metal1 656 -3300 656 -3300 5 vdd
rlabel metal1 629 -3300 629 -3300 5 vdd
rlabel metal1 648 -3497 648 -3497 1 gnd
rlabel metal1 1042 -2998 1042 -2998 1 gnd
rlabel metal1 1042 -2902 1042 -2902 5 vdd
rlabel metal1 999 -3029 999 -3029 1 gnd
rlabel metal1 1007 -2832 1007 -2832 5 vdd
rlabel metal1 980 -2832 980 -2832 5 vdd
rlabel metal1 1041 -2715 1041 -2715 1 gnd
rlabel metal1 1041 -2619 1041 -2619 5 vdd
rlabel metal1 998 -2746 998 -2746 1 gnd
rlabel metal1 1006 -2549 1006 -2549 5 vdd
rlabel metal1 979 -2549 979 -2549 5 vdd
rlabel metal1 708 -3733 708 -3733 1 gnd
rlabel metal1 708 -3637 708 -3637 5 vdd
rlabel metal1 665 -3764 665 -3764 1 gnd
rlabel metal1 673 -3567 673 -3567 5 vdd
rlabel metal1 646 -3567 646 -3567 5 vdd
rlabel metal1 696 -3982 696 -3982 1 gnd
rlabel metal1 696 -3886 696 -3886 5 vdd
rlabel metal1 661 -3816 661 -3816 5 vdd
rlabel metal1 634 -3816 634 -3816 5 vdd
rlabel metal1 653 -4013 653 -4013 1 gnd
rlabel metal1 1372 -3400 1372 -3400 1 gnd
rlabel metal1 1372 -3304 1372 -3304 5 vdd
rlabel metal1 1329 -3431 1329 -3431 1 gnd
rlabel metal1 1337 -3234 1337 -3234 5 vdd
rlabel metal1 1310 -3234 1310 -3234 5 vdd
rlabel metal1 1032 -3532 1032 -3532 1 gnd
rlabel metal1 1032 -3436 1032 -3436 5 vdd
rlabel metal1 997 -3366 997 -3366 5 vdd
rlabel metal1 970 -3366 970 -3366 5 vdd
rlabel metal1 989 -3563 989 -3563 1 gnd
rlabel metal1 1813 -2804 1813 -2804 5 vdd
rlabel metal1 1798 -3047 1798 -3047 1 gnd
rlabel metal1 1831 -3047 1831 -3047 1 gnd
rlabel metal1 1862 -2941 1862 -2941 5 vdd
rlabel metal1 1862 -3037 1862 -3037 1 gnd
rlabel metal1 861 1594 861 1594 7 vdd
rlabel metal1 765 1594 765 1594 3 gnd
rlabel metal1 861 1645 861 1645 7 vdd
rlabel metal1 765 1645 765 1645 3 gnd
rlabel metal1 913 1587 913 1587 1 gnd
rlabel metal1 913 1683 913 1683 5 vdd
rlabel metal1 1240 1532 1240 1532 1 gnd
rlabel metal1 1240 1628 1240 1628 5 vdd
rlabel metal1 1197 1501 1197 1501 1 gnd
rlabel metal1 1205 1698 1205 1698 5 vdd
rlabel metal1 1178 1698 1178 1698 5 vdd
rlabel metal1 1118 1477 1118 1477 1 gnd
rlabel metal1 1118 1573 1118 1573 5 vdd
rlabel metal1 1087 1467 1087 1467 1 gnd
rlabel metal1 1054 1467 1054 1467 1 gnd
rlabel metal1 1069 1710 1069 1710 5 vdd
rlabel metal1 1004 1571 1004 1571 1 gnd
rlabel metal1 1004 1667 1004 1667 5 vdd
rlabel metal1 3052 1640 3052 1640 5 vdd
rlabel metal1 3052 1544 3052 1544 1 gnd
rlabel metal1 3117 1683 3117 1683 5 vdd
rlabel metal1 3102 1440 3102 1440 1 gnd
rlabel metal1 3135 1440 3135 1440 1 gnd
rlabel metal1 3166 1546 3166 1546 5 vdd
rlabel metal1 3166 1450 3166 1450 1 gnd
rlabel metal1 3226 1671 3226 1671 5 vdd
rlabel metal1 3253 1671 3253 1671 5 vdd
rlabel metal1 3245 1474 3245 1474 1 gnd
rlabel metal1 3288 1601 3288 1601 5 vdd
rlabel metal1 3288 1505 3288 1505 1 gnd
rlabel metal1 2961 1656 2961 1656 5 vdd
rlabel metal1 2961 1560 2961 1560 1 gnd
rlabel metal1 2813 1618 2813 1618 3 gnd
rlabel metal1 2909 1618 2909 1618 7 vdd
rlabel metal1 2813 1567 2813 1567 3 gnd
rlabel metal1 2909 1567 2909 1567 7 vdd
rlabel metal1 3773 407 3773 407 5 vdd
rlabel metal1 3773 242 3773 242 1 gnd
rlabel metal1 3825 407 3825 407 5 vdd
rlabel metal1 3825 242 3825 242 1 gnd
rlabel metal1 3877 242 3877 242 1 gnd
rlabel metal1 3877 407 3877 407 5 vdd
rlabel metal1 3929 242 3929 242 1 gnd
rlabel metal1 3929 407 3929 407 5 vdd
rlabel metal1 3746 317 3746 317 1 d
rlabel metal1 4005 313 4005 313 1 gnd
rlabel metal1 4006 415 4006 415 5 vdd
rlabel metal1 3973 313 3973 313 1 gnd
rlabel metal1 3974 415 3974 415 5 vdd
rlabel metal1 3752 228 3752 228 1 clk
rlabel metal1 3777 348 3777 348 1 d1
rlabel metal1 3799 318 3799 318 1 a
rlabel metal1 3829 349 3829 349 1 d2
rlabel metal1 3851 317 3851 317 1 q1
rlabel metal1 3881 281 3881 281 1 d3
rlabel metal1 3904 316 3904 316 1 b
rlabel metal1 3933 280 3933 280 1 d4
rlabel metal1 3952 349 3952 349 1 qmid
rlabel metal1 3987 349 3987 349 1 qnot
rlabel metal1 4017 350 4017 350 7 q
rlabel metal1 -1522 410 -1522 410 5 vdd
rlabel metal1 -1522 245 -1522 245 1 gnd
rlabel metal1 -1470 410 -1470 410 5 vdd
rlabel metal1 -1470 245 -1470 245 1 gnd
rlabel metal1 -1418 245 -1418 245 1 gnd
rlabel metal1 -1418 410 -1418 410 5 vdd
rlabel metal1 -1366 245 -1366 245 1 gnd
rlabel metal1 -1366 410 -1366 410 5 vdd
rlabel metal1 -1290 316 -1290 316 1 gnd
rlabel metal1 -1289 418 -1289 418 5 vdd
rlabel metal1 -1322 316 -1322 316 1 gnd
rlabel metal1 -1321 418 -1321 418 5 vdd
rlabel metal1 -1543 231 -1543 231 1 clk
rlabel metal1 -396 9 -396 9 5 vdd
rlabel metal1 -396 -156 -396 -156 1 gnd
rlabel metal1 -344 9 -344 9 5 vdd
rlabel metal1 -344 -156 -344 -156 1 gnd
rlabel metal1 -292 -156 -292 -156 1 gnd
rlabel metal1 -292 9 -292 9 5 vdd
rlabel metal1 -240 -156 -240 -156 1 gnd
rlabel metal1 -240 9 -240 9 5 vdd
rlabel metal1 -164 -85 -164 -85 1 gnd
rlabel metal1 -163 17 -163 17 5 vdd
rlabel metal1 -196 -85 -196 -85 1 gnd
rlabel metal1 -195 17 -195 17 5 vdd
rlabel metal1 -417 -170 -417 -170 1 clk
rlabel metal1 -400 -246 -400 -246 5 vdd
rlabel metal1 -400 -411 -400 -411 1 gnd
rlabel metal1 -348 -246 -348 -246 5 vdd
rlabel metal1 -348 -411 -348 -411 1 gnd
rlabel metal1 -296 -411 -296 -411 1 gnd
rlabel metal1 -296 -246 -296 -246 5 vdd
rlabel metal1 -244 -411 -244 -411 1 gnd
rlabel metal1 -244 -246 -244 -246 5 vdd
rlabel metal1 -168 -340 -168 -340 1 gnd
rlabel metal1 -167 -238 -167 -238 5 vdd
rlabel metal1 -200 -340 -200 -340 1 gnd
rlabel metal1 -199 -238 -199 -238 5 vdd
rlabel metal1 -421 -425 -421 -425 1 clk
rlabel metal1 -303 -828 -303 -828 5 vdd
rlabel metal1 -303 -993 -303 -993 1 gnd
rlabel metal1 -251 -828 -251 -828 5 vdd
rlabel metal1 -251 -993 -251 -993 1 gnd
rlabel metal1 -199 -993 -199 -993 1 gnd
rlabel metal1 -199 -828 -199 -828 5 vdd
rlabel metal1 -147 -993 -147 -993 1 gnd
rlabel metal1 -147 -828 -147 -828 5 vdd
rlabel metal1 -71 -922 -71 -922 1 gnd
rlabel metal1 -70 -820 -70 -820 5 vdd
rlabel metal1 -103 -922 -103 -922 1 gnd
rlabel metal1 -102 -820 -102 -820 5 vdd
rlabel metal1 -324 -1007 -324 -1007 1 clk
rlabel metal1 -343 -1230 -343 -1230 1 clk
rlabel metal1 -121 -1043 -121 -1043 5 vdd
rlabel metal1 -122 -1145 -122 -1145 1 gnd
rlabel metal1 -89 -1043 -89 -1043 5 vdd
rlabel metal1 -90 -1145 -90 -1145 1 gnd
rlabel metal1 -166 -1051 -166 -1051 5 vdd
rlabel metal1 -166 -1216 -166 -1216 1 gnd
rlabel metal1 -218 -1051 -218 -1051 5 vdd
rlabel metal1 -218 -1216 -218 -1216 1 gnd
rlabel metal1 -270 -1216 -270 -1216 1 gnd
rlabel metal1 -270 -1051 -270 -1051 5 vdd
rlabel metal1 -322 -1216 -322 -1216 1 gnd
rlabel metal1 -322 -1051 -322 -1051 5 vdd
rlabel metal1 -343 -1568 -343 -1568 1 clk
rlabel metal1 -121 -1381 -121 -1381 5 vdd
rlabel metal1 -122 -1483 -122 -1483 1 gnd
rlabel metal1 -89 -1381 -89 -1381 5 vdd
rlabel metal1 -90 -1483 -90 -1483 1 gnd
rlabel metal1 -166 -1389 -166 -1389 5 vdd
rlabel metal1 -166 -1554 -166 -1554 1 gnd
rlabel metal1 -218 -1389 -218 -1389 5 vdd
rlabel metal1 -218 -1554 -218 -1554 1 gnd
rlabel metal1 -270 -1554 -270 -1554 1 gnd
rlabel metal1 -270 -1389 -270 -1389 5 vdd
rlabel metal1 -322 -1554 -322 -1554 1 gnd
rlabel metal1 -322 -1389 -322 -1389 5 vdd
rlabel metal1 -337 -1726 -337 -1726 5 vdd
rlabel metal1 -337 -1891 -337 -1891 1 gnd
rlabel metal1 -285 -1726 -285 -1726 5 vdd
rlabel metal1 -285 -1891 -285 -1891 1 gnd
rlabel metal1 -233 -1891 -233 -1891 1 gnd
rlabel metal1 -233 -1726 -233 -1726 5 vdd
rlabel metal1 -181 -1891 -181 -1891 1 gnd
rlabel metal1 -181 -1726 -181 -1726 5 vdd
rlabel metal1 -105 -1820 -105 -1820 1 gnd
rlabel metal1 -104 -1718 -104 -1718 5 vdd
rlabel metal1 -137 -1820 -137 -1820 1 gnd
rlabel metal1 -136 -1718 -136 -1718 5 vdd
rlabel metal1 -358 -1905 -358 -1905 1 clk
rlabel metal1 -358 -2512 -358 -2512 1 clk
rlabel metal1 -136 -2325 -136 -2325 5 vdd
rlabel metal1 -137 -2427 -137 -2427 1 gnd
rlabel metal1 -104 -2325 -104 -2325 5 vdd
rlabel metal1 -105 -2427 -105 -2427 1 gnd
rlabel metal1 -181 -2333 -181 -2333 5 vdd
rlabel metal1 -181 -2498 -181 -2498 1 gnd
rlabel metal1 -233 -2333 -233 -2333 5 vdd
rlabel metal1 -233 -2498 -233 -2498 1 gnd
rlabel metal1 -285 -2498 -285 -2498 1 gnd
rlabel metal1 -285 -2333 -285 -2333 5 vdd
rlabel metal1 -337 -2498 -337 -2498 1 gnd
rlabel metal1 -337 -2333 -337 -2333 5 vdd
rlabel metal1 -337 -2603 -337 -2603 5 vdd
rlabel metal1 -337 -2768 -337 -2768 1 gnd
rlabel metal1 -285 -2603 -285 -2603 5 vdd
rlabel metal1 -285 -2768 -285 -2768 1 gnd
rlabel metal1 -233 -2768 -233 -2768 1 gnd
rlabel metal1 -233 -2603 -233 -2603 5 vdd
rlabel metal1 -181 -2768 -181 -2768 1 gnd
rlabel metal1 -181 -2603 -181 -2603 5 vdd
rlabel metal1 -105 -2697 -105 -2697 1 gnd
rlabel metal1 -104 -2595 -104 -2595 5 vdd
rlabel metal1 -137 -2697 -137 -2697 1 gnd
rlabel metal1 -136 -2595 -136 -2595 5 vdd
rlabel metal1 -358 -2782 -358 -2782 1 clk
rlabel metal1 1425 104 1425 104 5 vdd
rlabel metal1 1425 -61 1425 -61 1 gnd
rlabel metal1 1477 104 1477 104 5 vdd
rlabel metal1 1477 -61 1477 -61 1 gnd
rlabel metal1 1529 -61 1529 -61 1 gnd
rlabel metal1 1529 104 1529 104 5 vdd
rlabel metal1 1581 -61 1581 -61 1 gnd
rlabel metal1 1581 104 1581 104 5 vdd
rlabel metal1 1657 10 1657 10 1 gnd
rlabel metal1 1658 112 1658 112 5 vdd
rlabel metal1 1625 10 1625 10 1 gnd
rlabel metal1 1626 112 1626 112 5 vdd
rlabel metal1 1404 -75 1404 -75 1 clk
rlabel metal1 1440 -172 1440 -172 5 vdd
rlabel metal1 1440 -337 1440 -337 1 gnd
rlabel metal1 1492 -172 1492 -172 5 vdd
rlabel metal1 1492 -337 1492 -337 1 gnd
rlabel metal1 1544 -337 1544 -337 1 gnd
rlabel metal1 1544 -172 1544 -172 5 vdd
rlabel metal1 1596 -337 1596 -337 1 gnd
rlabel metal1 1596 -172 1596 -172 5 vdd
rlabel metal1 1672 -266 1672 -266 1 gnd
rlabel metal1 1673 -164 1673 -164 5 vdd
rlabel metal1 1640 -266 1640 -266 1 gnd
rlabel metal1 1641 -164 1641 -164 5 vdd
rlabel metal1 1419 -351 1419 -351 1 clk
rlabel metal1 1824 -845 1824 -845 5 vdd
rlabel metal1 1824 -1010 1824 -1010 1 gnd
rlabel metal1 1876 -845 1876 -845 5 vdd
rlabel metal1 1876 -1010 1876 -1010 1 gnd
rlabel metal1 1928 -1010 1928 -1010 1 gnd
rlabel metal1 1928 -845 1928 -845 5 vdd
rlabel metal1 1980 -1010 1980 -1010 1 gnd
rlabel metal1 1980 -845 1980 -845 5 vdd
rlabel metal1 2056 -939 2056 -939 1 gnd
rlabel metal1 2057 -837 2057 -837 5 vdd
rlabel metal1 2024 -939 2024 -939 1 gnd
rlabel metal1 2025 -837 2025 -837 5 vdd
rlabel metal1 1803 -1024 1803 -1024 1 clk
rlabel metal1 2013 -1595 2013 -1595 5 vdd
rlabel metal1 2013 -1760 2013 -1760 1 gnd
rlabel metal1 2065 -1595 2065 -1595 5 vdd
rlabel metal1 2065 -1760 2065 -1760 1 gnd
rlabel metal1 2117 -1760 2117 -1760 1 gnd
rlabel metal1 2117 -1595 2117 -1595 5 vdd
rlabel metal1 2169 -1760 2169 -1760 1 gnd
rlabel metal1 2169 -1595 2169 -1595 5 vdd
rlabel metal1 2245 -1689 2245 -1689 1 gnd
rlabel metal1 2246 -1587 2246 -1587 5 vdd
rlabel metal1 2213 -1689 2213 -1689 1 gnd
rlabel metal1 2214 -1587 2214 -1587 5 vdd
rlabel metal1 1992 -1774 1992 -1774 1 clk
rlabel metal1 2087 -2837 2087 -2837 5 vdd
rlabel metal1 2087 -3002 2087 -3002 1 gnd
rlabel metal1 2139 -2837 2139 -2837 5 vdd
rlabel metal1 2139 -3002 2139 -3002 1 gnd
rlabel metal1 2191 -3002 2191 -3002 1 gnd
rlabel metal1 2191 -2837 2191 -2837 5 vdd
rlabel metal1 2243 -3002 2243 -3002 1 gnd
rlabel metal1 2243 -2837 2243 -2837 5 vdd
rlabel metal1 2319 -2931 2319 -2931 1 gnd
rlabel metal1 2320 -2829 2320 -2829 5 vdd
rlabel metal1 2287 -2931 2287 -2931 1 gnd
rlabel metal1 2288 -2829 2288 -2829 5 vdd
rlabel metal1 2066 -3016 2066 -3016 1 clk
rlabel metal1 -423 -82 -423 -82 1 a0
rlabel metal1 -426 -343 -426 -343 1 b0
rlabel metal1 -330 -922 -330 -922 1 a1
rlabel metal1 -349 -1149 -349 -1149 1 b1
rlabel metal1 -348 -1488 -348 -1488 1 a2
rlabel metal1 -363 -1824 -363 -1824 1 b2
rlabel metal1 -363 -2430 -363 -2430 1 a3
rlabel metal1 -364 -2700 -364 -2700 1 b3
rlabel metal1 1670 46 1671 47 1 s0
rlabel metal1 1686 -231 1687 -230 1 s1
rlabel metal1 2070 -902 2071 -901 1 s2
rlabel metal1 2257 -1654 2258 -1653 1 s3
rlabel metal1 2334 -2895 2335 -2894 1 cout
rlabel metal1 1894 -3003 1894 -3003 1 C4
<< end >>
